module file_handler();
  


endmodule;