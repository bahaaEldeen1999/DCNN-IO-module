
// 	Thu May  6 06:57:58 2021
//	vlsi
//	localhost.localdomain

module DMA (address, data, read_signal, write_signal, dataout, clk, RST, doneRead, 
    doneWrite);

output [15:0] dataout;
output doneRead;
output doneWrite;
input RST;
input [15:0] address;
input clk;
input [15:0] data;
input read_signal;
input write_signal;
wire \mem[10][15] ;
wire \mem[10][14] ;
wire \mem[10][13] ;
wire \mem[10][12] ;
wire \mem[10][11] ;
wire \mem[10][10] ;
wire \mem[10][9] ;
wire \mem[10][8] ;
wire \mem[10][7] ;
wire \mem[10][6] ;
wire \mem[10][5] ;
wire \mem[10][4] ;
wire \mem[10][3] ;
wire \mem[10][2] ;
wire \mem[10][1] ;
wire \mem[10][0] ;
wire \mem[9][15] ;
wire \mem[9][14] ;
wire \mem[9][13] ;
wire \mem[9][12] ;
wire \mem[9][11] ;
wire \mem[9][10] ;
wire \mem[9][9] ;
wire \mem[9][8] ;
wire \mem[9][7] ;
wire \mem[9][6] ;
wire \mem[9][5] ;
wire \mem[9][4] ;
wire \mem[9][3] ;
wire \mem[9][2] ;
wire \mem[9][1] ;
wire \mem[9][0] ;
wire \mem[8][15] ;
wire \mem[8][14] ;
wire \mem[8][13] ;
wire \mem[8][12] ;
wire \mem[8][11] ;
wire \mem[8][10] ;
wire \mem[8][9] ;
wire \mem[8][8] ;
wire \mem[8][7] ;
wire \mem[8][6] ;
wire \mem[8][5] ;
wire \mem[8][4] ;
wire \mem[8][3] ;
wire \mem[8][2] ;
wire \mem[8][1] ;
wire \mem[8][0] ;
wire \mem[7][15] ;
wire \mem[7][14] ;
wire \mem[7][13] ;
wire \mem[7][12] ;
wire \mem[7][11] ;
wire \mem[7][10] ;
wire \mem[7][9] ;
wire \mem[7][8] ;
wire \mem[7][7] ;
wire \mem[7][6] ;
wire \mem[7][5] ;
wire \mem[7][4] ;
wire \mem[7][3] ;
wire \mem[7][2] ;
wire \mem[7][1] ;
wire \mem[7][0] ;
wire \mem[6][15] ;
wire \mem[6][14] ;
wire \mem[6][13] ;
wire \mem[6][12] ;
wire \mem[6][11] ;
wire \mem[6][10] ;
wire \mem[6][9] ;
wire \mem[6][8] ;
wire \mem[6][7] ;
wire \mem[6][6] ;
wire \mem[6][5] ;
wire \mem[6][4] ;
wire \mem[6][3] ;
wire \mem[6][2] ;
wire \mem[6][1] ;
wire \mem[6][0] ;
wire \mem[5][15] ;
wire \mem[5][14] ;
wire \mem[5][13] ;
wire \mem[5][12] ;
wire \mem[5][11] ;
wire \mem[5][10] ;
wire \mem[5][9] ;
wire \mem[5][8] ;
wire \mem[5][7] ;
wire \mem[5][6] ;
wire \mem[5][5] ;
wire \mem[5][4] ;
wire \mem[5][3] ;
wire \mem[5][2] ;
wire \mem[5][1] ;
wire \mem[5][0] ;
wire \mem[4][15] ;
wire \mem[4][14] ;
wire \mem[4][13] ;
wire \mem[4][12] ;
wire \mem[4][11] ;
wire \mem[4][10] ;
wire \mem[4][9] ;
wire \mem[4][8] ;
wire \mem[4][7] ;
wire \mem[4][6] ;
wire \mem[4][5] ;
wire \mem[4][4] ;
wire \mem[4][3] ;
wire \mem[4][2] ;
wire \mem[4][1] ;
wire \mem[4][0] ;
wire \mem[1][15] ;
wire \mem[1][14] ;
wire \mem[1][13] ;
wire \mem[1][12] ;
wire \mem[1][11] ;
wire \mem[1][10] ;
wire \mem[1][9] ;
wire \mem[1][8] ;
wire \mem[1][7] ;
wire \mem[1][6] ;
wire \mem[1][5] ;
wire \mem[1][4] ;
wire \mem[1][3] ;
wire \mem[1][2] ;
wire \mem[1][1] ;
wire \mem[1][0] ;
wire n_0_13;
wire n_0_191_0;
wire n_0_191_1;
wire n_0_191_2;
wire n_0_31;
wire n_0_192_0;
wire n_0_192_1;
wire n_0_192_2;
wire n_0_10;
wire n_0_100_0;
wire n_0_100_1;
wire n_0_12;
wire n_0_117_0;
wire n_0_117_1;
wire n_0_14;
wire n_0_151_0;
wire n_0_151_1;
wire n_0_32;
wire \mem[3][15] ;
wire \mem[3][14] ;
wire \mem[3][13] ;
wire \mem[3][12] ;
wire \mem[3][11] ;
wire \mem[3][10] ;
wire \mem[3][9] ;
wire \mem[3][8] ;
wire \mem[3][7] ;
wire \mem[3][6] ;
wire \mem[3][5] ;
wire \mem[3][4] ;
wire \mem[3][3] ;
wire \mem[3][2] ;
wire \mem[3][1] ;
wire \mem[3][0] ;
wire \mem[2][15] ;
wire \mem[2][14] ;
wire \mem[2][13] ;
wire \mem[2][12] ;
wire \mem[2][11] ;
wire \mem[2][10] ;
wire \mem[2][9] ;
wire \mem[2][8] ;
wire \mem[2][7] ;
wire \mem[2][6] ;
wire \mem[2][5] ;
wire \mem[2][4] ;
wire \mem[2][3] ;
wire \mem[2][2] ;
wire \mem[2][1] ;
wire \mem[2][0] ;
wire \mem[0][15] ;
wire \mem[0][14] ;
wire \mem[0][13] ;
wire \mem[0][12] ;
wire \mem[0][11] ;
wire \mem[0][10] ;
wire \mem[0][9] ;
wire \mem[0][8] ;
wire \mem[0][7] ;
wire \mem[0][6] ;
wire \mem[0][5] ;
wire \mem[0][4] ;
wire \mem[0][3] ;
wire \mem[0][2] ;
wire \mem[0][1] ;
wire \mem[0][0] ;
wire n_0_0_0;
wire n_0_0_1;
wire n_0_0_2;
wire n_0_0_3;
wire n_0_0_4;
wire n_0_0_5;
wire n_0_0_6;
wire n_0_0_7;
wire n_0_0_8;
wire n_0_0_9;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_0_14;
wire n_0_0_15;
wire n_0_0_16;
wire n_0_0_17;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_0_21;
wire n_0_0_22;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_0_28;
wire n_0_0_29;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_0_32;
wire n_0_0_33;
wire n_0_0_34;
wire n_0_48;
wire n_0_5_20;
wire n_0_69;
wire n_0_5_0;
wire n_0_5_1;
wire n_0_5_2;
wire n_0_5_3;
wire n_0_5_4;
wire n_0_5_5;
wire n_0_5_6;
wire n_0_5_7;
wire n_0_5_8;
wire n_0_5_9;
wire n_0_5_10;
wire n_0_5_11;
wire n_0_5_12;
wire n_0_5_13;
wire n_0_5_14;
wire n_0_5_15;
wire n_0_5_16;
wire n_0_5_17;
wire n_0_5_18;
wire n_0_5_19;
wire n_0_5_21;
wire n_0_5_22;
wire n_0_5_23;
wire n_0_5_24;
wire n_0_5_25;
wire n_0_5_26;
wire n_0_5_27;
wire n_0_5_28;
wire n_0_5_29;
wire n_0_5_30;
wire n_0_5_31;
wire n_0_5_32;
wire n_0_5_33;
wire n_0_5_34;
wire n_0_5_35;
wire n_0_5_36;
wire n_0_8_0;
wire n_0_8_2;
wire n_0_8_3;
wire n_0_8_4;
wire n_0_8_5;
wire n_0_8_6;
wire n_0_8_7;
wire n_0_8_1;
wire n_0_8_9;
wire n_0_8_10;
wire n_0_8_11;
wire n_0_8_12;
wire n_0_8_13;
wire n_0_8_14;
wire n_0_8_15;
wire n_0_8_16;
wire n_0_8_17;
wire n_0_8_18;
wire n_0_8_19;
wire n_0_8_20;
wire n_0_8_21;
wire n_0_8_22;
wire n_0_8_23;
wire n_0_8_24;
wire n_0_8_25;
wire n_0_8_26;
wire n_0_8_27;
wire n_0_8_28;
wire n_0_8_8;
wire n_0_8_29;
wire n_0_8_30;
wire n_0_8_31;
wire n_0_8_32;
wire n_0_8_33;
wire n_0_8_34;
wire n_0_70;
wire n_0_15;
wire n_0_9_0;
wire n_0_9_1;
wire n_0_9_2;
wire n_0_9_3;
wire n_0_9_4;
wire n_0_9_5;
wire n_0_9_6;
wire n_0_9_7;
wire n_0_9_8;
wire n_0_9_9;
wire n_0_9_10;
wire n_0_9_11;
wire n_0_9_12;
wire n_0_9_13;
wire n_0_9_14;
wire n_0_9_15;
wire n_0_9_16;
wire n_0_9_17;
wire n_0_9_18;
wire n_0_9_19;
wire n_0_9_20;
wire n_0_9_21;
wire n_0_9_22;
wire n_0_9_23;
wire n_0_9_24;
wire n_0_9_25;
wire n_0_9_26;
wire n_0_9_27;
wire n_0_9_28;
wire n_0_9_29;
wire n_0_9_30;
wire n_0_9_31;
wire n_0_9_32;
wire n_0_9_33;
wire n_0_9_34;
wire n_0_16;
wire n_0_10_0;
wire n_0_10_1;
wire n_0_10_2;
wire n_0_10_3;
wire n_0_10_4;
wire n_0_10_5;
wire n_0_10_6;
wire n_0_10_7;
wire n_0_10_8;
wire n_0_10_9;
wire n_0_10_10;
wire n_0_10_11;
wire n_0_10_12;
wire n_0_10_13;
wire n_0_10_14;
wire n_0_10_15;
wire n_0_10_16;
wire n_0_10_17;
wire n_0_10_18;
wire n_0_10_19;
wire n_0_10_20;
wire n_0_10_21;
wire n_0_10_22;
wire n_0_10_23;
wire n_0_10_24;
wire n_0_10_25;
wire n_0_10_26;
wire n_0_10_27;
wire n_0_10_28;
wire n_0_10_29;
wire n_0_10_30;
wire n_0_10_31;
wire n_0_10_32;
wire n_0_10_33;
wire n_0_10_34;
wire n_0_17_0;
wire n_0_17_1;
wire n_0_17_2;
wire n_0_17_3;
wire n_0_17_4;
wire n_0_17_5;
wire n_0_17_6;
wire n_0_17_7;
wire n_0_17_8;
wire n_0_17_9;
wire n_0_17_10;
wire n_0_17_11;
wire n_0_17_12;
wire n_0_17_13;
wire n_0_17_14;
wire n_0_17_15;
wire n_0_17_16;
wire n_0_17_17;
wire n_0_17_18;
wire n_0_17_19;
wire n_0_17_20;
wire n_0_17_21;
wire n_0_17_22;
wire n_0_17_23;
wire n_0_17_24;
wire n_0_17;
wire n_0_17_25;
wire n_0_17_26;
wire n_0_17_27;
wire n_0_17_28;
wire n_0_17_29;
wire n_0_17_30;
wire n_0_17_31;
wire n_0_17_32;
wire n_0_17_33;
wire n_0_34_0;
wire n_0_34_1;
wire n_0_34_2;
wire n_0_34_3;
wire n_0_34_4;
wire n_0_34_5;
wire n_0_34_6;
wire n_0_34_7;
wire n_0_34_8;
wire n_0_34_9;
wire n_0_34_10;
wire n_0_34_11;
wire n_0_34_12;
wire n_0_34_13;
wire n_0_34_14;
wire n_0_34_15;
wire n_0_34_16;
wire n_0_34_17;
wire n_0_34_18;
wire n_0_34_19;
wire n_0_34_20;
wire n_0_34_21;
wire n_0_34_22;
wire n_0_34_23;
wire n_0_34_24;
wire n_0_18;
wire n_0_34_25;
wire n_0_34_26;
wire n_0_34_27;
wire n_0_34_28;
wire n_0_34_29;
wire n_0_34_30;
wire n_0_34_31;
wire n_0_34_32;
wire n_0_34_33;
wire n_0_51_0;
wire n_0_51_1;
wire n_0_51_2;
wire n_0_51_3;
wire n_0_51_4;
wire n_0_51_5;
wire n_0_51_6;
wire n_0_51_7;
wire n_0_51_8;
wire n_0_51_9;
wire n_0_51_10;
wire n_0_51_11;
wire n_0_51_12;
wire n_0_51_13;
wire n_0_51_14;
wire n_0_51_15;
wire n_0_51_16;
wire n_0_51_17;
wire n_0_51_18;
wire n_0_51_19;
wire n_0_51_20;
wire n_0_51_21;
wire n_0_51_22;
wire n_0_51_23;
wire n_0_51_24;
wire n_0_51_25;
wire n_0_51_26;
wire n_0_51_27;
wire n_0_51_28;
wire n_0_51_29;
wire n_0_51_30;
wire n_0_51_31;
wire n_0_51_32;
wire n_0_51_33;
wire n_0_51_34;
wire n_0_19;
wire n_0_20;
wire n_0_68_0;
wire n_0_68_1;
wire n_0_68_2;
wire n_0_68_3;
wire n_0_68_4;
wire n_0_68_5;
wire n_0_68_6;
wire n_0_68_7;
wire n_0_68_8;
wire n_0_68_9;
wire n_0_68_10;
wire n_0_68_11;
wire n_0_68_12;
wire n_0_68_13;
wire n_0_68_14;
wire n_0_68_15;
wire n_0_68_16;
wire n_0_68_17;
wire n_0_68_18;
wire n_0_68_19;
wire n_0_68_20;
wire n_0_68_21;
wire n_0_68_22;
wire n_0_68_23;
wire n_0_68_24;
wire n_0_68_25;
wire n_0_68_26;
wire n_0_21;
wire n_0_85_0;
wire n_0_85_1;
wire n_0_85_2;
wire n_0_85_3;
wire n_0_85_4;
wire n_0_85_5;
wire n_0_85_6;
wire n_0_85_7;
wire n_0_85_8;
wire n_0_85_9;
wire n_0_85_10;
wire n_0_85_11;
wire n_0_85_12;
wire n_0_85_13;
wire n_0_85_14;
wire n_0_85_15;
wire n_0_85_16;
wire n_0_85_17;
wire n_0_85_18;
wire n_0_85_19;
wire n_0_85_20;
wire n_0_85_21;
wire n_0_85_22;
wire n_0_85_23;
wire n_0_85_24;
wire n_0_85_25;
wire n_0_85_26;
wire n_0_85_27;
wire n_0_85_28;
wire n_0_85_29;
wire n_0_85_30;
wire n_0_22;
wire n_0_102_0;
wire n_0_102_1;
wire n_0_102_2;
wire n_0_102_3;
wire n_0_102_4;
wire n_0_102_5;
wire n_0_102_6;
wire n_0_102_7;
wire n_0_102_8;
wire n_0_102_9;
wire n_0_102_10;
wire n_0_102_11;
wire n_0_102_12;
wire n_0_102_13;
wire n_0_102_14;
wire n_0_102_15;
wire n_0_102_16;
wire n_0_102_17;
wire n_0_102_18;
wire n_0_102_19;
wire n_0_102_20;
wire n_0_102_21;
wire n_0_102_22;
wire n_0_102_23;
wire n_0_102_24;
wire n_0_102_25;
wire n_0_102_26;
wire n_0_102_27;
wire n_0_102_28;
wire n_0_102_29;
wire n_0_102_30;
wire n_0_119_0;
wire n_0_119_1;
wire n_0_119_2;
wire n_0_119_3;
wire n_0_119_4;
wire n_0_119_5;
wire n_0_119_6;
wire n_0_119_7;
wire n_0_119_8;
wire n_0_119_9;
wire n_0_119_10;
wire n_0_119_11;
wire n_0_119_12;
wire n_0_119_13;
wire n_0_119_14;
wire n_0_119_15;
wire n_0_119_16;
wire n_0_119_17;
wire n_0_119_18;
wire n_0_119_19;
wire n_0_119_20;
wire n_0_119_21;
wire n_0_119_22;
wire n_0_119_23;
wire n_0_119_24;
wire n_0_119_25;
wire n_0_119_26;
wire n_0_119_27;
wire n_0_119_28;
wire n_0_119_29;
wire n_0_119_30;
wire n_0_119_31;
wire n_0_119_32;
wire n_0_119_33;
wire n_0_119_34;
wire n_0_119_35;
wire n_0_23;
wire n_0_24;
wire n_0_136_0;
wire n_0_136_1;
wire n_0_136_2;
wire n_0_136_3;
wire n_0_136_4;
wire n_0_136_5;
wire n_0_136_6;
wire n_0_136_7;
wire n_0_136_8;
wire n_0_136_9;
wire n_0_136_10;
wire n_0_136_11;
wire n_0_136_12;
wire n_0_136_13;
wire n_0_136_14;
wire n_0_136_15;
wire n_0_136_16;
wire n_0_136_17;
wire n_0_136_18;
wire n_0_136_19;
wire n_0_136_20;
wire n_0_136_21;
wire n_0_136_22;
wire n_0_136_23;
wire n_0_136_24;
wire n_0_136_25;
wire n_0_136_26;
wire n_0_136_27;
wire n_0_136_28;
wire n_0_136_29;
wire n_0_136_30;
wire n_0_153_0;
wire n_0_153_1;
wire n_0_153_2;
wire n_0_153_3;
wire n_0_153_4;
wire n_0_153_5;
wire n_0_153_6;
wire n_0_153_7;
wire n_0_153_8;
wire n_0_153_9;
wire n_0_153_10;
wire n_0_153_11;
wire n_0_153_12;
wire n_0_153_13;
wire n_0_153_14;
wire n_0_153_15;
wire n_0_153_16;
wire n_0_153_17;
wire n_0_153_18;
wire n_0_153_19;
wire n_0_153_20;
wire n_0_153_21;
wire n_0_153_22;
wire n_0_153_23;
wire n_0_153_24;
wire n_0_153_25;
wire n_0_153_26;
wire n_0_153_27;
wire n_0_153_28;
wire n_0_153_29;
wire n_0_153_30;
wire n_0_153_31;
wire n_0_153_32;
wire n_0_153_33;
wire n_0_153_34;
wire n_0_153_35;
wire n_0_25;
wire n_0_170_0;
wire n_0_170_1;
wire n_0_170_2;
wire n_0_170_3;
wire n_0_170_4;
wire n_0_170_5;
wire n_0_170_6;
wire n_0_170_7;
wire n_0_170_8;
wire n_0_170_9;
wire n_0_170_10;
wire n_0_170_11;
wire n_0_170_12;
wire n_0_170_13;
wire n_0_170_14;
wire n_0_170_15;
wire n_0_170_16;
wire n_0_170_17;
wire n_0_170_18;
wire n_0_170_19;
wire n_0_170_20;
wire n_0_170_21;
wire n_0_170_22;
wire n_0_170_23;
wire n_0_170_24;
wire n_0_170_25;
wire n_0_170_26;
wire n_0_170_27;
wire n_0_170_28;
wire n_0_170_29;
wire n_0_170_30;
wire n_0_170_31;
wire n_0_170_32;
wire n_0_170_33;
wire n_0_170_34;
wire n_0_170_35;
wire n_0_26;
wire n_0_18_0;
wire n_0_18_1;
wire n_0_18_2;
wire n_0_18_3;
wire n_0_18_4;
wire n_0_18_5;
wire n_0_18_6;
wire n_0_18_7;
wire n_0_18_8;
wire n_0_18_9;
wire n_0_18_10;
wire n_0_18_11;
wire n_0_18_12;
wire n_0_18_13;
wire n_0_18_14;
wire n_0_18_15;
wire n_0_18_16;
wire n_0_18_17;
wire n_0_18_18;
wire n_0_18_19;
wire n_0_18_20;
wire n_0_18_21;
wire n_0_18_22;
wire n_0_18_23;
wire n_0_18_24;
wire n_0_18_25;
wire n_0_18_26;
wire n_0_18_27;
wire n_0_18_28;
wire n_0_18_29;
wire n_0_18_30;
wire n_0_18_31;
wire n_0_18_32;
wire n_0_18_33;
wire n_0_18_34;
wire n_0_18_35;
wire n_0_18_36;
wire n_0_27;
wire n_0_35_0;
wire n_0_35_1;
wire n_0_35_2;
wire n_0_35_3;
wire n_0_35_4;
wire n_0_35_5;
wire n_0_35_6;
wire n_0_35_7;
wire n_0_35_8;
wire n_0_35_9;
wire n_0_35_10;
wire n_0_35_11;
wire n_0_35_12;
wire n_0_35_13;
wire n_0_35_14;
wire n_0_35_15;
wire n_0_35_16;
wire n_0_35_17;
wire n_0_35_18;
wire n_0_35_19;
wire n_0_35_20;
wire n_0_35_21;
wire n_0_35_22;
wire n_0_35_23;
wire n_0_35_24;
wire n_0_28;
wire n_0_35_25;
wire n_0_35_26;
wire n_0_35_27;
wire n_0_35_28;
wire n_0_35_29;
wire n_0_35_30;
wire n_0_35_31;
wire n_0_35_32;
wire n_0_35_33;
wire n_0_52_0;
wire n_0_52_1;
wire n_0_52_2;
wire n_0_52_3;
wire n_0_52_4;
wire n_0_52_5;
wire n_0_52_6;
wire n_0_52_7;
wire n_0_52_8;
wire n_0_52_9;
wire n_0_52_10;
wire n_0_52_11;
wire n_0_52_12;
wire n_0_52_13;
wire n_0_52_14;
wire n_0_52_15;
wire n_0_52_16;
wire n_0_52_17;
wire n_0_52_18;
wire n_0_52_19;
wire n_0_52_20;
wire n_0_52_21;
wire n_0_52_22;
wire n_0_52_23;
wire n_0_52_24;
wire n_0_29;
wire n_0_52_25;
wire n_0_52_26;
wire n_0_52_27;
wire n_0_52_28;
wire n_0_52_29;
wire n_0_52_30;
wire n_0_52_31;
wire n_0_52_32;
wire n_0_52_33;
wire n_0_69_0;
wire n_0_69_1;
wire n_0_69_2;
wire n_0_69_3;
wire n_0_69_4;
wire n_0_69_5;
wire n_0_69_6;
wire n_0_69_7;
wire n_0_69_8;
wire n_0_69_9;
wire n_0_69_10;
wire n_0_69_11;
wire n_0_69_12;
wire n_0_69_13;
wire n_0_69_14;
wire n_0_69_15;
wire n_0_69_16;
wire n_0_69_17;
wire n_0_69_18;
wire n_0_69_19;
wire n_0_69_20;
wire n_0_69_21;
wire n_0_69_22;
wire n_0_69_23;
wire n_0_69_24;
wire n_0_69_25;
wire n_0_69_26;
wire n_0_69_27;
wire n_0_69_28;
wire n_0_69_29;
wire n_0_69_30;
wire n_0_69_31;
wire n_0_69_32;
wire n_0_69_33;
wire n_0_69_34;
wire n_0_30;
wire n_0_33;
wire n_0_86_0;
wire n_0_86_1;
wire n_0_86_2;
wire n_0_86_3;
wire n_0_86_4;
wire n_0_86_5;
wire n_0_86_6;
wire n_0_86_7;
wire n_0_86_8;
wire n_0_86_9;
wire n_0_86_10;
wire n_0_86_11;
wire n_0_86_12;
wire n_0_86_13;
wire n_0_86_14;
wire n_0_86_15;
wire n_0_86_16;
wire n_0_86_17;
wire n_0_86_18;
wire n_0_86_19;
wire n_0_86_20;
wire n_0_86_21;
wire n_0_86_22;
wire n_0_86_23;
wire n_0_86_24;
wire n_0_86_25;
wire n_0_86_26;
wire n_0_34;
wire n_0_103_0;
wire n_0_103_1;
wire n_0_103_2;
wire n_0_103_3;
wire n_0_103_4;
wire n_0_103_5;
wire n_0_103_6;
wire n_0_103_7;
wire n_0_103_8;
wire n_0_103_9;
wire n_0_103_10;
wire n_0_103_11;
wire n_0_103_12;
wire n_0_103_13;
wire n_0_103_14;
wire n_0_103_15;
wire n_0_103_16;
wire n_0_103_17;
wire n_0_103_18;
wire n_0_103_19;
wire n_0_103_20;
wire n_0_103_21;
wire n_0_103_22;
wire n_0_103_23;
wire n_0_103_24;
wire n_0_103_25;
wire n_0_103_26;
wire n_0_103_27;
wire n_0_103_28;
wire n_0_103_29;
wire n_0_103_30;
wire n_0_35;
wire n_0_120_0;
wire n_0_120_1;
wire n_0_120_2;
wire n_0_120_3;
wire n_0_120_4;
wire n_0_120_5;
wire n_0_120_6;
wire n_0_120_7;
wire n_0_120_8;
wire n_0_120_9;
wire n_0_120_10;
wire n_0_120_11;
wire n_0_120_12;
wire n_0_120_13;
wire n_0_120_14;
wire n_0_120_15;
wire n_0_120_16;
wire n_0_120_17;
wire n_0_120_18;
wire n_0_120_19;
wire n_0_120_20;
wire n_0_120_21;
wire n_0_120_22;
wire n_0_120_23;
wire n_0_120_24;
wire n_0_120_25;
wire n_0_120_26;
wire n_0_120_27;
wire n_0_120_28;
wire n_0_120_29;
wire n_0_120_30;
wire n_0_137_0;
wire n_0_137_1;
wire n_0_137_2;
wire n_0_137_3;
wire n_0_137_4;
wire n_0_137_5;
wire n_0_137_6;
wire n_0_137_7;
wire n_0_137_8;
wire n_0_137_9;
wire n_0_137_10;
wire n_0_137_11;
wire n_0_137_12;
wire n_0_137_13;
wire n_0_137_14;
wire n_0_137_15;
wire n_0_137_16;
wire n_0_137_17;
wire n_0_137_18;
wire n_0_137_19;
wire n_0_137_20;
wire n_0_137_21;
wire n_0_137_22;
wire n_0_137_23;
wire n_0_137_24;
wire n_0_137_25;
wire n_0_137_26;
wire n_0_137_27;
wire n_0_137_28;
wire n_0_137_29;
wire n_0_137_30;
wire n_0_137_31;
wire n_0_137_32;
wire n_0_137_33;
wire n_0_137_34;
wire n_0_137_35;
wire n_0_36;
wire n_0_37;
wire n_0_154_0;
wire n_0_154_1;
wire n_0_154_2;
wire n_0_154_3;
wire n_0_154_4;
wire n_0_154_5;
wire n_0_154_6;
wire n_0_154_7;
wire n_0_154_8;
wire n_0_154_9;
wire n_0_154_10;
wire n_0_154_11;
wire n_0_154_12;
wire n_0_154_13;
wire n_0_154_14;
wire n_0_154_15;
wire n_0_154_16;
wire n_0_154_17;
wire n_0_154_18;
wire n_0_154_19;
wire n_0_154_20;
wire n_0_154_21;
wire n_0_154_22;
wire n_0_154_23;
wire n_0_154_24;
wire n_0_154_25;
wire n_0_154_26;
wire n_0_154_27;
wire n_0_154_28;
wire n_0_154_29;
wire n_0_154_30;
wire n_0_171_0;
wire n_0_171_1;
wire n_0_171_2;
wire n_0_171_3;
wire n_0_171_4;
wire n_0_171_5;
wire n_0_171_6;
wire n_0_171_7;
wire n_0_171_8;
wire n_0_171_9;
wire n_0_171_10;
wire n_0_171_11;
wire n_0_171_12;
wire n_0_171_13;
wire n_0_171_14;
wire n_0_171_15;
wire n_0_171_16;
wire n_0_171_17;
wire n_0_171_18;
wire n_0_171_19;
wire n_0_171_20;
wire n_0_171_21;
wire n_0_171_22;
wire n_0_171_23;
wire n_0_171_24;
wire n_0_171_25;
wire n_0_171_26;
wire n_0_171_27;
wire n_0_171_28;
wire n_0_171_29;
wire n_0_171_30;
wire n_0_171_31;
wire n_0_171_32;
wire n_0_171_33;
wire n_0_171_34;
wire n_0_171_35;
wire n_0_38;
wire n_0_33_0;
wire n_0_33_1;
wire n_0_33_2;
wire n_0_33_3;
wire n_0_33_4;
wire n_0_33_5;
wire n_0_33_6;
wire n_0_33_7;
wire n_0_33_8;
wire n_0_33_9;
wire n_0_33_10;
wire n_0_33_11;
wire n_0_33_12;
wire n_0_33_13;
wire n_0_33_14;
wire n_0_33_15;
wire n_0_33_16;
wire n_0_33_17;
wire n_0_33_18;
wire n_0_33_19;
wire n_0_33_20;
wire n_0_33_21;
wire n_0_33_22;
wire n_0_33_23;
wire n_0_33_24;
wire n_0_33_25;
wire n_0_33_26;
wire n_0_33_27;
wire n_0_33_28;
wire n_0_33_29;
wire n_0_33_30;
wire n_0_33_31;
wire n_0_33_32;
wire n_0_33_33;
wire n_0_33_34;
wire n_0_33_35;
wire n_0_39;
wire n_0_19_0;
wire n_0_19_1;
wire n_0_19_2;
wire n_0_19_3;
wire n_0_19_4;
wire n_0_19_5;
wire n_0_19_6;
wire n_0_19_7;
wire n_0_19_8;
wire n_0_19_9;
wire n_0_19_10;
wire n_0_19_11;
wire n_0_19_12;
wire n_0_19_13;
wire n_0_19_14;
wire n_0_19_15;
wire n_0_19_16;
wire n_0_19_17;
wire n_0_19_18;
wire n_0_19_19;
wire n_0_19_20;
wire n_0_19_21;
wire n_0_19_22;
wire n_0_19_23;
wire n_0_19_24;
wire n_0_19_25;
wire n_0_19_26;
wire n_0_19_27;
wire n_0_19_28;
wire n_0_19_29;
wire n_0_19_30;
wire n_0_19_31;
wire n_0_19_32;
wire n_0_19_33;
wire n_0_19_34;
wire n_0_19_35;
wire n_0_19_36;
wire n_0_40;
wire n_0_36_0;
wire n_0_36_1;
wire n_0_36_2;
wire n_0_36_3;
wire n_0_36_4;
wire n_0_36_5;
wire n_0_36_6;
wire n_0_36_7;
wire n_0_36_8;
wire n_0_36_9;
wire n_0_36_10;
wire n_0_36_11;
wire n_0_36_12;
wire n_0_36_13;
wire n_0_36_14;
wire n_0_36_15;
wire n_0_36_16;
wire n_0_36_17;
wire n_0_36_18;
wire n_0_36_19;
wire n_0_36_20;
wire n_0_36_21;
wire n_0_36_22;
wire n_0_36_23;
wire n_0_36_24;
wire n_0_41;
wire n_0_36_25;
wire n_0_36_26;
wire n_0_36_27;
wire n_0_36_28;
wire n_0_36_29;
wire n_0_36_30;
wire n_0_36_31;
wire n_0_36_32;
wire n_0_36_33;
wire n_0_53_0;
wire n_0_53_1;
wire n_0_53_2;
wire n_0_53_3;
wire n_0_53_4;
wire n_0_53_5;
wire n_0_53_6;
wire n_0_53_7;
wire n_0_53_8;
wire n_0_53_9;
wire n_0_53_10;
wire n_0_53_11;
wire n_0_53_12;
wire n_0_53_13;
wire n_0_53_14;
wire n_0_53_15;
wire n_0_53_16;
wire n_0_53_17;
wire n_0_53_18;
wire n_0_53_19;
wire n_0_53_20;
wire n_0_53_21;
wire n_0_53_22;
wire n_0_53_23;
wire n_0_53_24;
wire n_0_42;
wire n_0_53_25;
wire n_0_53_26;
wire n_0_53_27;
wire n_0_53_28;
wire n_0_53_29;
wire n_0_53_30;
wire n_0_53_31;
wire n_0_53_32;
wire n_0_53_33;
wire n_0_70_0;
wire n_0_70_1;
wire n_0_70_2;
wire n_0_70_3;
wire n_0_70_4;
wire n_0_70_5;
wire n_0_70_6;
wire n_0_70_7;
wire n_0_70_8;
wire n_0_70_9;
wire n_0_70_10;
wire n_0_70_11;
wire n_0_70_12;
wire n_0_70_13;
wire n_0_70_14;
wire n_0_70_15;
wire n_0_70_16;
wire n_0_70_17;
wire n_0_70_18;
wire n_0_70_19;
wire n_0_70_20;
wire n_0_70_21;
wire n_0_70_22;
wire n_0_70_23;
wire n_0_70_24;
wire n_0_70_25;
wire n_0_70_26;
wire n_0_70_27;
wire n_0_70_28;
wire n_0_70_29;
wire n_0_70_30;
wire n_0_70_31;
wire n_0_70_32;
wire n_0_70_33;
wire n_0_70_34;
wire n_0_43;
wire n_0_44;
wire n_0_87_0;
wire n_0_87_1;
wire n_0_87_2;
wire n_0_87_3;
wire n_0_87_4;
wire n_0_87_5;
wire n_0_87_6;
wire n_0_87_7;
wire n_0_87_8;
wire n_0_87_9;
wire n_0_87_10;
wire n_0_87_11;
wire n_0_87_12;
wire n_0_87_13;
wire n_0_87_14;
wire n_0_87_15;
wire n_0_87_16;
wire n_0_87_17;
wire n_0_87_18;
wire n_0_87_19;
wire n_0_87_20;
wire n_0_87_21;
wire n_0_87_22;
wire n_0_87_23;
wire n_0_87_24;
wire n_0_87_25;
wire n_0_87_26;
wire n_0_45;
wire n_0_104_0;
wire n_0_104_1;
wire n_0_104_2;
wire n_0_104_3;
wire n_0_104_4;
wire n_0_104_5;
wire n_0_104_6;
wire n_0_104_7;
wire n_0_104_8;
wire n_0_104_9;
wire n_0_104_10;
wire n_0_104_11;
wire n_0_104_12;
wire n_0_104_13;
wire n_0_104_14;
wire n_0_104_15;
wire n_0_104_16;
wire n_0_104_17;
wire n_0_104_18;
wire n_0_104_19;
wire n_0_104_20;
wire n_0_104_21;
wire n_0_104_22;
wire n_0_104_23;
wire n_0_104_24;
wire n_0_104_25;
wire n_0_104_26;
wire n_0_104_27;
wire n_0_104_28;
wire n_0_104_29;
wire n_0_104_30;
wire n_0_46;
wire n_0_121_0;
wire n_0_121_1;
wire n_0_121_2;
wire n_0_121_3;
wire n_0_121_4;
wire n_0_121_5;
wire n_0_121_6;
wire n_0_121_7;
wire n_0_121_8;
wire n_0_121_9;
wire n_0_121_10;
wire n_0_121_11;
wire n_0_121_12;
wire n_0_121_13;
wire n_0_121_14;
wire n_0_121_15;
wire n_0_121_16;
wire n_0_121_17;
wire n_0_121_18;
wire n_0_121_19;
wire n_0_121_20;
wire n_0_121_21;
wire n_0_121_22;
wire n_0_121_23;
wire n_0_121_24;
wire n_0_121_25;
wire n_0_121_26;
wire n_0_121_27;
wire n_0_121_28;
wire n_0_121_29;
wire n_0_121_30;
wire n_0_138_0;
wire n_0_138_1;
wire n_0_138_2;
wire n_0_138_3;
wire n_0_138_4;
wire n_0_138_5;
wire n_0_138_6;
wire n_0_138_7;
wire n_0_138_8;
wire n_0_138_9;
wire n_0_138_10;
wire n_0_138_11;
wire n_0_138_12;
wire n_0_138_13;
wire n_0_138_14;
wire n_0_138_15;
wire n_0_138_16;
wire n_0_138_17;
wire n_0_138_18;
wire n_0_138_19;
wire n_0_138_20;
wire n_0_138_21;
wire n_0_138_22;
wire n_0_138_23;
wire n_0_138_24;
wire n_0_138_25;
wire n_0_138_26;
wire n_0_138_27;
wire n_0_138_28;
wire n_0_138_29;
wire n_0_138_30;
wire n_0_138_31;
wire n_0_138_32;
wire n_0_138_33;
wire n_0_138_34;
wire n_0_138_35;
wire n_0_47;
wire n_0_50;
wire n_0_155_0;
wire n_0_155_1;
wire n_0_155_2;
wire n_0_155_3;
wire n_0_155_4;
wire n_0_155_5;
wire n_0_155_6;
wire n_0_155_7;
wire n_0_155_8;
wire n_0_155_9;
wire n_0_155_10;
wire n_0_155_11;
wire n_0_155_12;
wire n_0_155_13;
wire n_0_155_14;
wire n_0_155_15;
wire n_0_155_16;
wire n_0_155_17;
wire n_0_155_18;
wire n_0_155_19;
wire n_0_155_20;
wire n_0_155_21;
wire n_0_155_22;
wire n_0_155_23;
wire n_0_155_24;
wire n_0_155_25;
wire n_0_155_26;
wire n_0_155_27;
wire n_0_155_28;
wire n_0_155_29;
wire n_0_155_30;
wire n_0_172_0;
wire n_0_172_1;
wire n_0_172_2;
wire n_0_172_3;
wire n_0_172_4;
wire n_0_172_5;
wire n_0_172_6;
wire n_0_172_7;
wire n_0_172_8;
wire n_0_172_9;
wire n_0_172_10;
wire n_0_172_11;
wire n_0_172_12;
wire n_0_172_13;
wire n_0_172_14;
wire n_0_172_15;
wire n_0_172_16;
wire n_0_172_17;
wire n_0_172_18;
wire n_0_172_19;
wire n_0_172_20;
wire n_0_172_21;
wire n_0_172_22;
wire n_0_172_23;
wire n_0_172_24;
wire n_0_172_25;
wire n_0_172_26;
wire n_0_172_27;
wire n_0_172_28;
wire n_0_172_29;
wire n_0_172_30;
wire n_0_172_31;
wire n_0_172_32;
wire n_0_172_33;
wire n_0_172_34;
wire n_0_172_35;
wire n_0_51;
wire n_0_50_0;
wire n_0_50_1;
wire n_0_50_2;
wire n_0_50_3;
wire n_0_50_4;
wire n_0_50_5;
wire n_0_50_6;
wire n_0_50_7;
wire n_0_50_8;
wire n_0_50_9;
wire n_0_50_10;
wire n_0_50_11;
wire n_0_50_12;
wire n_0_50_13;
wire n_0_50_14;
wire n_0_50_15;
wire n_0_50_16;
wire n_0_50_17;
wire n_0_50_18;
wire n_0_50_19;
wire n_0_50_20;
wire n_0_50_21;
wire n_0_50_22;
wire n_0_50_23;
wire n_0_50_24;
wire n_0_50_25;
wire n_0_50_26;
wire n_0_50_27;
wire n_0_50_28;
wire n_0_50_29;
wire n_0_50_30;
wire n_0_50_31;
wire n_0_50_32;
wire n_0_50_33;
wire n_0_50_34;
wire n_0_50_35;
wire n_0_52;
wire n_0_20_0;
wire n_0_20_1;
wire n_0_20_2;
wire n_0_20_3;
wire n_0_20_4;
wire n_0_20_5;
wire n_0_20_6;
wire n_0_20_7;
wire n_0_20_8;
wire n_0_20_9;
wire n_0_20_10;
wire n_0_20_11;
wire n_0_20_12;
wire n_0_20_13;
wire n_0_20_14;
wire n_0_20_15;
wire n_0_20_16;
wire n_0_20_17;
wire n_0_20_18;
wire n_0_20_19;
wire n_0_20_20;
wire n_0_20_21;
wire n_0_20_22;
wire n_0_20_23;
wire n_0_20_24;
wire n_0_20_25;
wire n_0_20_26;
wire n_0_20_27;
wire n_0_20_28;
wire n_0_20_29;
wire n_0_20_30;
wire n_0_20_31;
wire n_0_20_32;
wire n_0_20_33;
wire n_0_20_34;
wire n_0_20_35;
wire n_0_20_36;
wire n_0_53;
wire n_0_37_0;
wire n_0_37_1;
wire n_0_37_2;
wire n_0_37_3;
wire n_0_37_4;
wire n_0_37_5;
wire n_0_37_6;
wire n_0_37_7;
wire n_0_37_8;
wire n_0_37_9;
wire n_0_37_10;
wire n_0_37_11;
wire n_0_37_12;
wire n_0_37_13;
wire n_0_37_14;
wire n_0_37_15;
wire n_0_37_16;
wire n_0_37_17;
wire n_0_37_18;
wire n_0_37_19;
wire n_0_37_20;
wire n_0_37_21;
wire n_0_37_22;
wire n_0_37_23;
wire n_0_37_24;
wire n_0_54;
wire n_0_37_25;
wire n_0_37_26;
wire n_0_37_27;
wire n_0_37_28;
wire n_0_37_29;
wire n_0_37_30;
wire n_0_37_31;
wire n_0_37_32;
wire n_0_37_33;
wire n_0_54_0;
wire n_0_54_1;
wire n_0_54_2;
wire n_0_54_3;
wire n_0_54_4;
wire n_0_54_5;
wire n_0_54_6;
wire n_0_54_7;
wire n_0_54_8;
wire n_0_54_9;
wire n_0_54_10;
wire n_0_54_11;
wire n_0_54_12;
wire n_0_54_13;
wire n_0_54_14;
wire n_0_54_15;
wire n_0_54_16;
wire n_0_54_17;
wire n_0_54_18;
wire n_0_54_19;
wire n_0_54_20;
wire n_0_54_21;
wire n_0_54_22;
wire n_0_54_23;
wire n_0_54_24;
wire n_0_55;
wire n_0_54_25;
wire n_0_54_26;
wire n_0_54_27;
wire n_0_54_28;
wire n_0_54_29;
wire n_0_54_30;
wire n_0_54_31;
wire n_0_54_32;
wire n_0_54_33;
wire n_0_71_0;
wire n_0_71_1;
wire n_0_71_2;
wire n_0_71_3;
wire n_0_71_4;
wire n_0_71_5;
wire n_0_71_6;
wire n_0_71_7;
wire n_0_71_8;
wire n_0_71_9;
wire n_0_71_10;
wire n_0_71_11;
wire n_0_71_12;
wire n_0_71_13;
wire n_0_71_14;
wire n_0_71_15;
wire n_0_71_16;
wire n_0_71_17;
wire n_0_71_18;
wire n_0_71_19;
wire n_0_71_20;
wire n_0_71_21;
wire n_0_71_22;
wire n_0_71_23;
wire n_0_71_24;
wire n_0_71_25;
wire n_0_71_26;
wire n_0_71_27;
wire n_0_71_28;
wire n_0_71_29;
wire n_0_71_30;
wire n_0_71_31;
wire n_0_71_32;
wire n_0_71_33;
wire n_0_71_34;
wire n_0_56;
wire n_0_57;
wire n_0_88_0;
wire n_0_88_1;
wire n_0_88_2;
wire n_0_88_3;
wire n_0_88_4;
wire n_0_88_5;
wire n_0_88_6;
wire n_0_88_7;
wire n_0_88_8;
wire n_0_88_9;
wire n_0_88_10;
wire n_0_88_11;
wire n_0_88_12;
wire n_0_88_13;
wire n_0_88_14;
wire n_0_88_15;
wire n_0_88_16;
wire n_0_88_17;
wire n_0_88_18;
wire n_0_88_19;
wire n_0_88_20;
wire n_0_88_21;
wire n_0_88_22;
wire n_0_88_23;
wire n_0_88_24;
wire n_0_88_25;
wire n_0_88_26;
wire n_0_58;
wire n_0_105_0;
wire n_0_105_1;
wire n_0_105_2;
wire n_0_105_3;
wire n_0_105_4;
wire n_0_105_5;
wire n_0_105_6;
wire n_0_105_7;
wire n_0_105_8;
wire n_0_105_9;
wire n_0_105_10;
wire n_0_105_11;
wire n_0_105_12;
wire n_0_105_13;
wire n_0_105_14;
wire n_0_105_15;
wire n_0_105_16;
wire n_0_105_17;
wire n_0_105_18;
wire n_0_105_19;
wire n_0_105_20;
wire n_0_105_21;
wire n_0_105_22;
wire n_0_105_23;
wire n_0_105_24;
wire n_0_105_25;
wire n_0_105_26;
wire n_0_105_27;
wire n_0_105_28;
wire n_0_105_29;
wire n_0_105_30;
wire n_0_59;
wire n_0_122_0;
wire n_0_122_1;
wire n_0_122_2;
wire n_0_122_3;
wire n_0_122_4;
wire n_0_122_5;
wire n_0_122_6;
wire n_0_122_7;
wire n_0_122_8;
wire n_0_122_9;
wire n_0_122_10;
wire n_0_122_11;
wire n_0_122_12;
wire n_0_122_13;
wire n_0_122_14;
wire n_0_122_15;
wire n_0_122_16;
wire n_0_122_17;
wire n_0_122_18;
wire n_0_122_19;
wire n_0_122_20;
wire n_0_122_21;
wire n_0_122_22;
wire n_0_122_23;
wire n_0_122_24;
wire n_0_122_25;
wire n_0_122_26;
wire n_0_122_27;
wire n_0_122_28;
wire n_0_122_29;
wire n_0_122_30;
wire n_0_139_0;
wire n_0_139_1;
wire n_0_139_2;
wire n_0_139_3;
wire n_0_139_4;
wire n_0_139_5;
wire n_0_139_6;
wire n_0_139_7;
wire n_0_139_8;
wire n_0_139_9;
wire n_0_139_10;
wire n_0_139_11;
wire n_0_139_12;
wire n_0_139_13;
wire n_0_139_14;
wire n_0_139_15;
wire n_0_139_16;
wire n_0_139_17;
wire n_0_139_18;
wire n_0_139_19;
wire n_0_139_20;
wire n_0_139_21;
wire n_0_139_22;
wire n_0_139_23;
wire n_0_139_24;
wire n_0_139_25;
wire n_0_139_26;
wire n_0_139_27;
wire n_0_139_28;
wire n_0_139_29;
wire n_0_139_30;
wire n_0_139_31;
wire n_0_139_32;
wire n_0_139_33;
wire n_0_139_34;
wire n_0_139_35;
wire n_0_60;
wire n_0_61;
wire n_0_156_0;
wire n_0_156_1;
wire n_0_156_2;
wire n_0_156_3;
wire n_0_156_4;
wire n_0_156_5;
wire n_0_156_6;
wire n_0_156_7;
wire n_0_156_8;
wire n_0_156_9;
wire n_0_156_10;
wire n_0_156_11;
wire n_0_156_12;
wire n_0_156_13;
wire n_0_156_14;
wire n_0_156_15;
wire n_0_156_16;
wire n_0_156_17;
wire n_0_156_18;
wire n_0_156_19;
wire n_0_156_20;
wire n_0_156_21;
wire n_0_156_22;
wire n_0_156_23;
wire n_0_156_24;
wire n_0_156_25;
wire n_0_156_26;
wire n_0_156_27;
wire n_0_156_28;
wire n_0_156_29;
wire n_0_156_30;
wire n_0_173_0;
wire n_0_173_1;
wire n_0_173_2;
wire n_0_173_3;
wire n_0_173_4;
wire n_0_173_5;
wire n_0_173_6;
wire n_0_173_7;
wire n_0_173_8;
wire n_0_173_9;
wire n_0_173_10;
wire n_0_173_11;
wire n_0_173_12;
wire n_0_173_13;
wire n_0_173_14;
wire n_0_173_15;
wire n_0_173_16;
wire n_0_173_17;
wire n_0_173_18;
wire n_0_173_19;
wire n_0_173_20;
wire n_0_173_21;
wire n_0_173_22;
wire n_0_173_23;
wire n_0_173_24;
wire n_0_173_25;
wire n_0_173_26;
wire n_0_173_27;
wire n_0_173_28;
wire n_0_173_29;
wire n_0_173_30;
wire n_0_173_31;
wire n_0_173_32;
wire n_0_173_33;
wire n_0_173_34;
wire n_0_173_35;
wire n_0_62;
wire n_0_67_0;
wire n_0_67_1;
wire n_0_67_2;
wire n_0_67_3;
wire n_0_67_4;
wire n_0_67_5;
wire n_0_67_6;
wire n_0_67_7;
wire n_0_67_8;
wire n_0_67_9;
wire n_0_67_10;
wire n_0_67_11;
wire n_0_67_12;
wire n_0_67_13;
wire n_0_67_14;
wire n_0_67_15;
wire n_0_67_16;
wire n_0_67_17;
wire n_0_67_18;
wire n_0_67_19;
wire n_0_67_20;
wire n_0_67_21;
wire n_0_67_22;
wire n_0_67_23;
wire n_0_67_24;
wire n_0_67_25;
wire n_0_67_26;
wire n_0_67_27;
wire n_0_67_28;
wire n_0_67_29;
wire n_0_67_30;
wire n_0_67_31;
wire n_0_67_32;
wire n_0_67_33;
wire n_0_67_34;
wire n_0_67_35;
wire n_0_63;
wire n_0_3_0;
wire n_0_3_1;
wire n_0_3_2;
wire n_0_3_3;
wire n_0_3_4;
wire n_0_3_5;
wire n_0_3_6;
wire n_0_3_7;
wire n_0_3_8;
wire n_0_3_9;
wire n_0_3_10;
wire n_0_3_11;
wire n_0_3_12;
wire n_0_3_13;
wire n_0_3_14;
wire n_0_3_15;
wire n_0_3_16;
wire n_0_3_17;
wire n_0_3_18;
wire n_0_3_19;
wire n_0_3_20;
wire n_0_3_21;
wire n_0_3_22;
wire n_0_3_23;
wire n_0_3_24;
wire n_0_3_25;
wire n_0_3_26;
wire n_0_3_27;
wire n_0_3_28;
wire n_0_3_29;
wire n_0_3_30;
wire n_0_3_31;
wire n_0_3_32;
wire n_0_3_33;
wire n_0_3_34;
wire n_0_3_35;
wire n_0_3_36;
wire n_0_64;
wire n_0_21_20;
wire n_0_71;
wire n_0_21_0;
wire n_0_21_1;
wire n_0_21_2;
wire n_0_21_3;
wire n_0_21_4;
wire n_0_21_5;
wire n_0_21_6;
wire n_0_21_7;
wire n_0_21_8;
wire n_0_21_9;
wire n_0_21_10;
wire n_0_21_11;
wire n_0_21_12;
wire n_0_21_13;
wire n_0_21_14;
wire n_0_21_15;
wire n_0_21_16;
wire n_0_21_17;
wire n_0_21_18;
wire n_0_21_19;
wire n_0_21_21;
wire n_0_21_22;
wire n_0_21_23;
wire n_0_21_24;
wire n_0_21_25;
wire n_0_21_26;
wire n_0_21_27;
wire n_0_21_28;
wire n_0_21_29;
wire n_0_21_30;
wire n_0_21_31;
wire n_0_21_32;
wire n_0_21_33;
wire n_0_21_34;
wire n_0_21_35;
wire n_0_21_36;
wire n_0_38_0;
wire n_0_38_1;
wire n_0_38_2;
wire n_0_38_3;
wire n_0_38_4;
wire n_0_38_5;
wire n_0_38_6;
wire n_0_38_7;
wire n_0_38_8;
wire n_0_38_9;
wire n_0_38_10;
wire n_0_38_11;
wire n_0_38_12;
wire n_0_38_13;
wire n_0_38_14;
wire n_0_38_15;
wire n_0_38_16;
wire n_0_38_17;
wire n_0_38_18;
wire n_0_38_19;
wire n_0_38_20;
wire n_0_38_21;
wire n_0_38_22;
wire n_0_38_23;
wire n_0_38_24;
wire n_0_75;
wire n_0_38_25;
wire n_0_38_26;
wire n_0_38_27;
wire n_0_38_28;
wire n_0_38_29;
wire n_0_38_30;
wire n_0_38_31;
wire n_0_38_32;
wire n_0_38_33;
wire n_0_55_0;
wire n_0_55_1;
wire n_0_55_2;
wire n_0_55_3;
wire n_0_55_4;
wire n_0_55_5;
wire n_0_55_6;
wire n_0_55_7;
wire n_0_55_8;
wire n_0_55_9;
wire n_0_55_10;
wire n_0_55_11;
wire n_0_55_12;
wire n_0_55_13;
wire n_0_55_14;
wire n_0_55_15;
wire n_0_55_16;
wire n_0_55_17;
wire n_0_55_18;
wire n_0_55_19;
wire n_0_55_20;
wire n_0_55_21;
wire n_0_55_22;
wire n_0_55_23;
wire n_0_55_24;
wire n_0_76;
wire n_0_55_25;
wire n_0_55_26;
wire n_0_55_27;
wire n_0_55_28;
wire n_0_55_29;
wire n_0_55_30;
wire n_0_55_31;
wire n_0_55_32;
wire n_0_55_33;
wire n_0_72_0;
wire n_0_72_1;
wire n_0_72_2;
wire n_0_72_3;
wire n_0_72_4;
wire n_0_72_5;
wire n_0_72_6;
wire n_0_72_7;
wire n_0_72_8;
wire n_0_72_9;
wire n_0_72_10;
wire n_0_72_11;
wire n_0_72_12;
wire n_0_72_13;
wire n_0_72_14;
wire n_0_72_15;
wire n_0_72_16;
wire n_0_72_17;
wire n_0_72_18;
wire n_0_72_19;
wire n_0_72_20;
wire n_0_72_21;
wire n_0_72_22;
wire n_0_72_23;
wire n_0_72_24;
wire n_0_72_25;
wire n_0_72_26;
wire n_0_72_27;
wire n_0_72_28;
wire n_0_72_29;
wire n_0_72_30;
wire n_0_72_31;
wire n_0_72_32;
wire n_0_72_33;
wire n_0_72_34;
wire n_0_77;
wire n_0_78;
wire n_0_89_0;
wire n_0_89_1;
wire n_0_89_2;
wire n_0_89_3;
wire n_0_89_4;
wire n_0_89_5;
wire n_0_89_6;
wire n_0_89_7;
wire n_0_89_8;
wire n_0_89_9;
wire n_0_89_10;
wire n_0_89_11;
wire n_0_89_12;
wire n_0_89_13;
wire n_0_89_14;
wire n_0_89_15;
wire n_0_89_16;
wire n_0_89_17;
wire n_0_89_18;
wire n_0_89_19;
wire n_0_89_20;
wire n_0_89_21;
wire n_0_89_22;
wire n_0_89_23;
wire n_0_89_24;
wire n_0_89_25;
wire n_0_89_26;
wire n_0_79;
wire n_0_106_0;
wire n_0_106_1;
wire n_0_106_2;
wire n_0_106_3;
wire n_0_106_4;
wire n_0_106_5;
wire n_0_106_6;
wire n_0_106_7;
wire n_0_106_8;
wire n_0_106_9;
wire n_0_106_10;
wire n_0_106_11;
wire n_0_106_12;
wire n_0_106_13;
wire n_0_106_14;
wire n_0_106_15;
wire n_0_106_16;
wire n_0_106_17;
wire n_0_106_18;
wire n_0_106_19;
wire n_0_106_20;
wire n_0_106_21;
wire n_0_106_22;
wire n_0_106_23;
wire n_0_106_24;
wire n_0_106_25;
wire n_0_106_26;
wire n_0_106_27;
wire n_0_106_28;
wire n_0_106_29;
wire n_0_106_30;
wire n_0_80;
wire n_0_123_0;
wire n_0_123_1;
wire n_0_123_2;
wire n_0_123_3;
wire n_0_123_4;
wire n_0_123_5;
wire n_0_123_6;
wire n_0_123_7;
wire n_0_123_8;
wire n_0_123_9;
wire n_0_123_10;
wire n_0_123_11;
wire n_0_123_12;
wire n_0_123_13;
wire n_0_123_14;
wire n_0_123_15;
wire n_0_123_16;
wire n_0_123_17;
wire n_0_123_18;
wire n_0_123_19;
wire n_0_123_20;
wire n_0_123_21;
wire n_0_123_22;
wire n_0_123_23;
wire n_0_123_24;
wire n_0_123_25;
wire n_0_123_26;
wire n_0_123_27;
wire n_0_123_28;
wire n_0_123_29;
wire n_0_123_30;
wire n_0_140_0;
wire n_0_140_1;
wire n_0_140_2;
wire n_0_140_3;
wire n_0_140_4;
wire n_0_140_5;
wire n_0_140_6;
wire n_0_140_7;
wire n_0_140_8;
wire n_0_140_9;
wire n_0_140_10;
wire n_0_140_11;
wire n_0_140_12;
wire n_0_140_13;
wire n_0_140_14;
wire n_0_140_15;
wire n_0_140_16;
wire n_0_140_17;
wire n_0_140_18;
wire n_0_140_19;
wire n_0_140_20;
wire n_0_140_21;
wire n_0_140_22;
wire n_0_140_23;
wire n_0_140_24;
wire n_0_140_25;
wire n_0_140_26;
wire n_0_140_27;
wire n_0_140_28;
wire n_0_140_29;
wire n_0_140_30;
wire n_0_140_31;
wire n_0_140_32;
wire n_0_140_33;
wire n_0_140_34;
wire n_0_140_35;
wire n_0_81;
wire n_0_82;
wire n_0_157_0;
wire n_0_157_1;
wire n_0_157_2;
wire n_0_157_3;
wire n_0_157_4;
wire n_0_157_5;
wire n_0_157_6;
wire n_0_157_7;
wire n_0_157_8;
wire n_0_157_9;
wire n_0_157_10;
wire n_0_157_11;
wire n_0_157_12;
wire n_0_157_13;
wire n_0_157_14;
wire n_0_157_15;
wire n_0_157_16;
wire n_0_157_17;
wire n_0_157_18;
wire n_0_157_19;
wire n_0_157_20;
wire n_0_157_21;
wire n_0_157_22;
wire n_0_157_23;
wire n_0_157_24;
wire n_0_157_25;
wire n_0_157_26;
wire n_0_157_27;
wire n_0_157_28;
wire n_0_157_29;
wire n_0_157_30;
wire n_0_174_0;
wire n_0_174_1;
wire n_0_174_2;
wire n_0_174_3;
wire n_0_174_4;
wire n_0_174_5;
wire n_0_174_6;
wire n_0_174_7;
wire n_0_174_8;
wire n_0_174_9;
wire n_0_174_10;
wire n_0_174_11;
wire n_0_174_12;
wire n_0_174_13;
wire n_0_174_14;
wire n_0_174_15;
wire n_0_174_16;
wire n_0_174_17;
wire n_0_174_18;
wire n_0_174_19;
wire n_0_174_20;
wire n_0_174_21;
wire n_0_174_22;
wire n_0_174_23;
wire n_0_174_24;
wire n_0_174_25;
wire n_0_174_26;
wire n_0_174_27;
wire n_0_174_28;
wire n_0_174_29;
wire n_0_174_30;
wire n_0_174_31;
wire n_0_174_32;
wire n_0_174_33;
wire n_0_174_34;
wire n_0_174_35;
wire n_0_83;
wire n_0_16_0;
wire n_0_16_1;
wire n_0_16_2;
wire n_0_16_3;
wire n_0_16_4;
wire n_0_16_5;
wire n_0_16_6;
wire n_0_16_7;
wire n_0_16_8;
wire n_0_16_9;
wire n_0_16_10;
wire n_0_16_11;
wire n_0_16_12;
wire n_0_16_13;
wire n_0_16_14;
wire n_0_16_15;
wire n_0_16_16;
wire n_0_16_17;
wire n_0_16_18;
wire n_0_16_19;
wire n_0_16_20;
wire n_0_16_21;
wire n_0_16_22;
wire n_0_16_23;
wire n_0_16_24;
wire n_0_16_25;
wire n_0_16_26;
wire n_0_16_27;
wire n_0_16_28;
wire n_0_16_29;
wire n_0_16_30;
wire n_0_16_31;
wire n_0_16_32;
wire n_0_16_33;
wire n_0_16_34;
wire n_0_16_35;
wire n_0_84;
wire n_0_22_0;
wire n_0_22_1;
wire n_0_22_2;
wire n_0_22_3;
wire n_0_22_4;
wire n_0_22_5;
wire n_0_22_6;
wire n_0_22_7;
wire n_0_22_8;
wire n_0_22_9;
wire n_0_22_10;
wire n_0_22_11;
wire n_0_22_12;
wire n_0_22_13;
wire n_0_22_14;
wire n_0_22_15;
wire n_0_22_16;
wire n_0_22_17;
wire n_0_22_18;
wire n_0_22_19;
wire n_0_22_20;
wire n_0_22_21;
wire n_0_22_22;
wire n_0_22_23;
wire n_0_22_24;
wire n_0_22_25;
wire n_0_22_26;
wire n_0_22_27;
wire n_0_22_28;
wire n_0_22_29;
wire n_0_22_30;
wire n_0_22_31;
wire n_0_22_32;
wire n_0_22_33;
wire n_0_22_34;
wire n_0_22_35;
wire n_0_22_36;
wire n_0_85;
wire n_0_39_0;
wire n_0_39_1;
wire n_0_39_2;
wire n_0_39_3;
wire n_0_39_4;
wire n_0_39_5;
wire n_0_39_6;
wire n_0_39_7;
wire n_0_39_8;
wire n_0_39_9;
wire n_0_39_10;
wire n_0_39_11;
wire n_0_39_12;
wire n_0_39_13;
wire n_0_39_14;
wire n_0_39_15;
wire n_0_39_16;
wire n_0_39_17;
wire n_0_39_18;
wire n_0_39_19;
wire n_0_39_20;
wire n_0_39_21;
wire n_0_39_22;
wire n_0_39_23;
wire n_0_39_24;
wire n_0_86;
wire n_0_39_25;
wire n_0_39_26;
wire n_0_39_27;
wire n_0_39_28;
wire n_0_39_29;
wire n_0_39_30;
wire n_0_39_31;
wire n_0_39_32;
wire n_0_39_33;
wire n_0_56_0;
wire n_0_56_1;
wire n_0_56_2;
wire n_0_56_3;
wire n_0_56_4;
wire n_0_56_5;
wire n_0_56_6;
wire n_0_56_7;
wire n_0_56_8;
wire n_0_56_9;
wire n_0_56_10;
wire n_0_56_11;
wire n_0_56_12;
wire n_0_56_13;
wire n_0_56_14;
wire n_0_56_15;
wire n_0_56_16;
wire n_0_56_17;
wire n_0_56_18;
wire n_0_56_19;
wire n_0_56_20;
wire n_0_56_21;
wire n_0_56_22;
wire n_0_56_23;
wire n_0_56_24;
wire n_0_87;
wire n_0_56_25;
wire n_0_56_26;
wire n_0_56_27;
wire n_0_56_28;
wire n_0_56_29;
wire n_0_56_30;
wire n_0_56_31;
wire n_0_56_32;
wire n_0_56_33;
wire n_0_73_0;
wire n_0_73_1;
wire n_0_73_2;
wire n_0_73_3;
wire n_0_73_4;
wire n_0_73_5;
wire n_0_73_6;
wire n_0_73_7;
wire n_0_73_8;
wire n_0_73_9;
wire n_0_73_10;
wire n_0_73_11;
wire n_0_73_12;
wire n_0_73_13;
wire n_0_73_14;
wire n_0_73_15;
wire n_0_73_16;
wire n_0_73_17;
wire n_0_73_18;
wire n_0_73_19;
wire n_0_73_20;
wire n_0_73_21;
wire n_0_73_22;
wire n_0_73_23;
wire n_0_73_24;
wire n_0_73_25;
wire n_0_73_26;
wire n_0_73_27;
wire n_0_73_28;
wire n_0_73_29;
wire n_0_73_30;
wire n_0_73_31;
wire n_0_73_32;
wire n_0_73_33;
wire n_0_73_34;
wire n_0_88;
wire n_0_89;
wire n_0_90_0;
wire n_0_90_1;
wire n_0_90_2;
wire n_0_90_3;
wire n_0_90_4;
wire n_0_90_5;
wire n_0_90_6;
wire n_0_90_7;
wire n_0_90_8;
wire n_0_90_9;
wire n_0_90_10;
wire n_0_90_11;
wire n_0_90_12;
wire n_0_90_13;
wire n_0_90_14;
wire n_0_90_15;
wire n_0_90_16;
wire n_0_90_17;
wire n_0_90_18;
wire n_0_90_19;
wire n_0_90_20;
wire n_0_90_21;
wire n_0_90_22;
wire n_0_90_23;
wire n_0_90_24;
wire n_0_90_25;
wire n_0_90_26;
wire n_0_90;
wire n_0_107_0;
wire n_0_107_1;
wire n_0_107_2;
wire n_0_107_3;
wire n_0_107_4;
wire n_0_107_5;
wire n_0_107_6;
wire n_0_107_7;
wire n_0_107_8;
wire n_0_107_9;
wire n_0_107_10;
wire n_0_107_11;
wire n_0_107_12;
wire n_0_107_13;
wire n_0_107_14;
wire n_0_107_15;
wire n_0_107_16;
wire n_0_107_17;
wire n_0_107_18;
wire n_0_107_19;
wire n_0_107_20;
wire n_0_107_21;
wire n_0_107_22;
wire n_0_107_23;
wire n_0_107_24;
wire n_0_107_25;
wire n_0_107_26;
wire n_0_107_27;
wire n_0_107_28;
wire n_0_107_29;
wire n_0_107_30;
wire n_0_91;
wire n_0_124_0;
wire n_0_124_1;
wire n_0_124_2;
wire n_0_124_3;
wire n_0_124_4;
wire n_0_124_5;
wire n_0_124_6;
wire n_0_124_7;
wire n_0_124_8;
wire n_0_124_9;
wire n_0_124_10;
wire n_0_124_11;
wire n_0_124_12;
wire n_0_124_13;
wire n_0_124_14;
wire n_0_124_15;
wire n_0_124_16;
wire n_0_124_17;
wire n_0_124_18;
wire n_0_124_19;
wire n_0_124_20;
wire n_0_124_21;
wire n_0_124_22;
wire n_0_124_23;
wire n_0_124_24;
wire n_0_124_25;
wire n_0_124_26;
wire n_0_124_27;
wire n_0_124_28;
wire n_0_124_29;
wire n_0_124_30;
wire n_0_141_0;
wire n_0_141_1;
wire n_0_141_2;
wire n_0_141_3;
wire n_0_141_4;
wire n_0_141_5;
wire n_0_141_6;
wire n_0_141_7;
wire n_0_141_8;
wire n_0_141_9;
wire n_0_141_10;
wire n_0_141_11;
wire n_0_141_12;
wire n_0_141_13;
wire n_0_141_14;
wire n_0_141_15;
wire n_0_141_16;
wire n_0_141_17;
wire n_0_141_18;
wire n_0_141_19;
wire n_0_141_20;
wire n_0_141_21;
wire n_0_141_22;
wire n_0_141_23;
wire n_0_141_24;
wire n_0_141_25;
wire n_0_141_26;
wire n_0_141_27;
wire n_0_141_28;
wire n_0_141_29;
wire n_0_141_30;
wire n_0_141_31;
wire n_0_141_32;
wire n_0_141_33;
wire n_0_141_34;
wire n_0_141_35;
wire n_0_92;
wire n_0_93;
wire n_0_158_0;
wire n_0_158_1;
wire n_0_158_2;
wire n_0_158_3;
wire n_0_158_4;
wire n_0_158_5;
wire n_0_158_6;
wire n_0_158_7;
wire n_0_158_8;
wire n_0_158_9;
wire n_0_158_10;
wire n_0_158_11;
wire n_0_158_12;
wire n_0_158_13;
wire n_0_158_14;
wire n_0_158_15;
wire n_0_158_16;
wire n_0_158_17;
wire n_0_158_18;
wire n_0_158_19;
wire n_0_158_20;
wire n_0_158_21;
wire n_0_158_22;
wire n_0_158_23;
wire n_0_158_24;
wire n_0_158_25;
wire n_0_158_26;
wire n_0_158_27;
wire n_0_158_28;
wire n_0_158_29;
wire n_0_158_30;
wire n_0_175_0;
wire n_0_175_1;
wire n_0_175_2;
wire n_0_175_3;
wire n_0_175_4;
wire n_0_175_5;
wire n_0_175_6;
wire n_0_175_7;
wire n_0_175_8;
wire n_0_175_9;
wire n_0_175_10;
wire n_0_175_11;
wire n_0_175_12;
wire n_0_175_13;
wire n_0_175_14;
wire n_0_175_15;
wire n_0_175_16;
wire n_0_175_17;
wire n_0_175_18;
wire n_0_175_19;
wire n_0_175_20;
wire n_0_175_21;
wire n_0_175_22;
wire n_0_175_23;
wire n_0_175_24;
wire n_0_175_25;
wire n_0_175_26;
wire n_0_175_27;
wire n_0_175_28;
wire n_0_175_29;
wire n_0_175_30;
wire n_0_175_31;
wire n_0_175_32;
wire n_0_175_33;
wire n_0_175_34;
wire n_0_175_35;
wire n_0_94;
wire n_0_101_0;
wire n_0_101_1;
wire n_0_101_2;
wire n_0_101_3;
wire n_0_101_4;
wire n_0_101_5;
wire n_0_101_6;
wire n_0_101_7;
wire n_0_101_8;
wire n_0_101_9;
wire n_0_101_10;
wire n_0_101_11;
wire n_0_101_12;
wire n_0_101_13;
wire n_0_101_14;
wire n_0_101_15;
wire n_0_101_16;
wire n_0_101_17;
wire n_0_101_18;
wire n_0_101_19;
wire n_0_101_20;
wire n_0_101_21;
wire n_0_101_22;
wire n_0_101_23;
wire n_0_101_24;
wire n_0_101_25;
wire n_0_101_26;
wire n_0_101_27;
wire n_0_101_28;
wire n_0_101_29;
wire n_0_101_30;
wire n_0_101_31;
wire n_0_101_32;
wire n_0_101_33;
wire n_0_101_34;
wire n_0_101_35;
wire n_0_95;
wire n_0_23_0;
wire n_0_23_1;
wire n_0_23_2;
wire n_0_23_3;
wire n_0_23_4;
wire n_0_23_5;
wire n_0_23_6;
wire n_0_23_7;
wire n_0_23_8;
wire n_0_23_9;
wire n_0_23_10;
wire n_0_23_11;
wire n_0_23_12;
wire n_0_23_13;
wire n_0_23_14;
wire n_0_23_15;
wire n_0_23_16;
wire n_0_23_17;
wire n_0_23_18;
wire n_0_23_19;
wire n_0_23_20;
wire n_0_23_21;
wire n_0_23_22;
wire n_0_23_23;
wire n_0_23_24;
wire n_0_23_25;
wire n_0_23_26;
wire n_0_23_27;
wire n_0_23_28;
wire n_0_23_29;
wire n_0_23_30;
wire n_0_23_31;
wire n_0_23_32;
wire n_0_23_33;
wire n_0_23_34;
wire n_0_23_35;
wire n_0_23_36;
wire n_0_96;
wire n_0_40_0;
wire n_0_40_1;
wire n_0_40_2;
wire n_0_40_3;
wire n_0_40_4;
wire n_0_40_5;
wire n_0_40_6;
wire n_0_40_7;
wire n_0_40_8;
wire n_0_40_9;
wire n_0_40_10;
wire n_0_40_11;
wire n_0_40_12;
wire n_0_40_13;
wire n_0_40_14;
wire n_0_40_15;
wire n_0_40_16;
wire n_0_40_17;
wire n_0_40_18;
wire n_0_40_19;
wire n_0_40_20;
wire n_0_40_21;
wire n_0_40_22;
wire n_0_40_23;
wire n_0_40_24;
wire n_0_97;
wire n_0_40_25;
wire n_0_40_26;
wire n_0_40_27;
wire n_0_40_28;
wire n_0_40_29;
wire n_0_40_30;
wire n_0_40_31;
wire n_0_40_32;
wire n_0_40_33;
wire n_0_57_0;
wire n_0_57_1;
wire n_0_57_2;
wire n_0_57_3;
wire n_0_57_4;
wire n_0_57_5;
wire n_0_57_6;
wire n_0_57_7;
wire n_0_57_8;
wire n_0_57_9;
wire n_0_57_10;
wire n_0_57_11;
wire n_0_57_12;
wire n_0_57_13;
wire n_0_57_14;
wire n_0_57_15;
wire n_0_57_16;
wire n_0_57_17;
wire n_0_57_18;
wire n_0_57_19;
wire n_0_57_20;
wire n_0_57_21;
wire n_0_57_22;
wire n_0_57_23;
wire n_0_57_24;
wire n_0_98;
wire n_0_57_25;
wire n_0_57_26;
wire n_0_57_27;
wire n_0_57_28;
wire n_0_57_29;
wire n_0_57_30;
wire n_0_57_31;
wire n_0_57_32;
wire n_0_57_33;
wire n_0_74_0;
wire n_0_74_1;
wire n_0_74_2;
wire n_0_74_3;
wire n_0_74_4;
wire n_0_74_5;
wire n_0_74_6;
wire n_0_74_7;
wire n_0_74_8;
wire n_0_74_9;
wire n_0_74_10;
wire n_0_74_11;
wire n_0_74_12;
wire n_0_74_13;
wire n_0_74_14;
wire n_0_74_15;
wire n_0_74_16;
wire n_0_74_17;
wire n_0_74_18;
wire n_0_74_19;
wire n_0_74_20;
wire n_0_74_21;
wire n_0_74_22;
wire n_0_74_23;
wire n_0_74_24;
wire n_0_74_25;
wire n_0_74_26;
wire n_0_74_27;
wire n_0_74_28;
wire n_0_74_29;
wire n_0_74_30;
wire n_0_74_31;
wire n_0_74_32;
wire n_0_74_33;
wire n_0_74_34;
wire n_0_101;
wire n_0_102;
wire n_0_91_0;
wire n_0_91_1;
wire n_0_91_2;
wire n_0_91_3;
wire n_0_91_4;
wire n_0_91_5;
wire n_0_91_6;
wire n_0_91_7;
wire n_0_91_8;
wire n_0_91_9;
wire n_0_91_10;
wire n_0_91_11;
wire n_0_91_12;
wire n_0_91_13;
wire n_0_91_14;
wire n_0_91_15;
wire n_0_91_16;
wire n_0_91_17;
wire n_0_91_18;
wire n_0_91_19;
wire n_0_91_20;
wire n_0_91_21;
wire n_0_91_22;
wire n_0_91_23;
wire n_0_91_24;
wire n_0_91_25;
wire n_0_91_26;
wire n_0_103;
wire n_0_108_0;
wire n_0_108_1;
wire n_0_108_2;
wire n_0_108_3;
wire n_0_108_4;
wire n_0_108_5;
wire n_0_108_6;
wire n_0_108_7;
wire n_0_108_8;
wire n_0_108_9;
wire n_0_108_10;
wire n_0_108_11;
wire n_0_108_12;
wire n_0_108_13;
wire n_0_108_14;
wire n_0_108_15;
wire n_0_108_16;
wire n_0_108_17;
wire n_0_108_18;
wire n_0_108_19;
wire n_0_108_20;
wire n_0_108_21;
wire n_0_108_22;
wire n_0_108_23;
wire n_0_108_24;
wire n_0_108_25;
wire n_0_108_26;
wire n_0_108_27;
wire n_0_108_28;
wire n_0_108_29;
wire n_0_108_30;
wire n_0_104;
wire n_0_125_0;
wire n_0_125_1;
wire n_0_125_2;
wire n_0_125_3;
wire n_0_125_4;
wire n_0_125_5;
wire n_0_125_6;
wire n_0_125_7;
wire n_0_125_8;
wire n_0_125_9;
wire n_0_125_10;
wire n_0_125_11;
wire n_0_125_12;
wire n_0_125_13;
wire n_0_125_14;
wire n_0_125_15;
wire n_0_125_16;
wire n_0_125_17;
wire n_0_125_18;
wire n_0_125_19;
wire n_0_125_20;
wire n_0_125_21;
wire n_0_125_22;
wire n_0_125_23;
wire n_0_125_24;
wire n_0_125_25;
wire n_0_125_26;
wire n_0_125_27;
wire n_0_125_28;
wire n_0_125_29;
wire n_0_125_30;
wire n_0_142_0;
wire n_0_142_1;
wire n_0_142_2;
wire n_0_142_3;
wire n_0_142_4;
wire n_0_142_5;
wire n_0_142_6;
wire n_0_142_7;
wire n_0_142_8;
wire n_0_142_9;
wire n_0_142_10;
wire n_0_142_11;
wire n_0_142_12;
wire n_0_142_13;
wire n_0_142_14;
wire n_0_142_15;
wire n_0_142_16;
wire n_0_142_17;
wire n_0_142_18;
wire n_0_142_19;
wire n_0_142_20;
wire n_0_142_21;
wire n_0_142_22;
wire n_0_142_23;
wire n_0_142_24;
wire n_0_142_25;
wire n_0_142_26;
wire n_0_142_27;
wire n_0_142_28;
wire n_0_142_29;
wire n_0_142_30;
wire n_0_142_31;
wire n_0_142_32;
wire n_0_142_33;
wire n_0_142_34;
wire n_0_142_35;
wire n_0_105;
wire n_0_106;
wire n_0_159_0;
wire n_0_159_1;
wire n_0_159_2;
wire n_0_159_3;
wire n_0_159_4;
wire n_0_159_5;
wire n_0_159_6;
wire n_0_159_7;
wire n_0_159_8;
wire n_0_159_9;
wire n_0_159_10;
wire n_0_159_11;
wire n_0_159_12;
wire n_0_159_13;
wire n_0_159_14;
wire n_0_159_15;
wire n_0_159_16;
wire n_0_159_17;
wire n_0_159_18;
wire n_0_159_19;
wire n_0_159_20;
wire n_0_159_21;
wire n_0_159_22;
wire n_0_159_23;
wire n_0_159_24;
wire n_0_159_25;
wire n_0_159_26;
wire n_0_159_27;
wire n_0_159_28;
wire n_0_159_29;
wire n_0_159_30;
wire n_0_176_0;
wire n_0_176_1;
wire n_0_176_2;
wire n_0_176_3;
wire n_0_176_4;
wire n_0_176_5;
wire n_0_176_6;
wire n_0_176_7;
wire n_0_176_8;
wire n_0_176_9;
wire n_0_176_10;
wire n_0_176_11;
wire n_0_176_12;
wire n_0_176_13;
wire n_0_176_14;
wire n_0_176_15;
wire n_0_176_16;
wire n_0_176_17;
wire n_0_176_18;
wire n_0_176_19;
wire n_0_176_20;
wire n_0_176_21;
wire n_0_176_22;
wire n_0_176_23;
wire n_0_176_24;
wire n_0_176_25;
wire n_0_176_26;
wire n_0_176_27;
wire n_0_176_28;
wire n_0_176_29;
wire n_0_176_30;
wire n_0_176_31;
wire n_0_176_32;
wire n_0_176_33;
wire n_0_176_34;
wire n_0_176_35;
wire n_0_107;
wire n_0_118_0;
wire n_0_118_1;
wire n_0_118_2;
wire n_0_118_3;
wire n_0_118_4;
wire n_0_118_5;
wire n_0_118_6;
wire n_0_118_7;
wire n_0_118_8;
wire n_0_118_9;
wire n_0_118_10;
wire n_0_118_11;
wire n_0_118_12;
wire n_0_118_13;
wire n_0_118_14;
wire n_0_118_15;
wire n_0_118_16;
wire n_0_118_17;
wire n_0_118_18;
wire n_0_118_19;
wire n_0_118_20;
wire n_0_118_21;
wire n_0_118_22;
wire n_0_118_23;
wire n_0_118_24;
wire n_0_118_25;
wire n_0_118_26;
wire n_0_118_27;
wire n_0_118_28;
wire n_0_118_29;
wire n_0_118_30;
wire n_0_118_31;
wire n_0_118_32;
wire n_0_118_33;
wire n_0_118_34;
wire n_0_118_35;
wire n_0_108;
wire n_0_24_0;
wire n_0_24_1;
wire n_0_24_2;
wire n_0_24_3;
wire n_0_24_4;
wire n_0_24_5;
wire n_0_24_6;
wire n_0_24_7;
wire n_0_24_8;
wire n_0_24_9;
wire n_0_24_10;
wire n_0_24_11;
wire n_0_24_12;
wire n_0_24_13;
wire n_0_24_14;
wire n_0_24_15;
wire n_0_24_16;
wire n_0_24_17;
wire n_0_24_18;
wire n_0_24_19;
wire n_0_24_20;
wire n_0_24_21;
wire n_0_24_22;
wire n_0_24_23;
wire n_0_24_24;
wire n_0_24_25;
wire n_0_24_26;
wire n_0_24_27;
wire n_0_24_28;
wire n_0_24_29;
wire n_0_24_30;
wire n_0_24_31;
wire n_0_24_32;
wire n_0_24_33;
wire n_0_24_34;
wire n_0_24_35;
wire n_0_24_36;
wire n_0_109;
wire n_0_41_0;
wire n_0_41_1;
wire n_0_41_2;
wire n_0_41_3;
wire n_0_41_4;
wire n_0_41_5;
wire n_0_41_6;
wire n_0_41_7;
wire n_0_41_8;
wire n_0_41_9;
wire n_0_41_10;
wire n_0_41_11;
wire n_0_41_12;
wire n_0_41_13;
wire n_0_41_14;
wire n_0_41_15;
wire n_0_41_16;
wire n_0_41_17;
wire n_0_41_18;
wire n_0_41_19;
wire n_0_41_20;
wire n_0_41_21;
wire n_0_41_22;
wire n_0_41_23;
wire n_0_41_24;
wire n_0_110;
wire n_0_41_25;
wire n_0_41_26;
wire n_0_41_27;
wire n_0_41_28;
wire n_0_41_29;
wire n_0_41_30;
wire n_0_41_31;
wire n_0_41_32;
wire n_0_41_33;
wire n_0_58_0;
wire n_0_58_1;
wire n_0_58_2;
wire n_0_58_3;
wire n_0_58_4;
wire n_0_58_5;
wire n_0_58_6;
wire n_0_58_7;
wire n_0_58_8;
wire n_0_58_9;
wire n_0_58_10;
wire n_0_58_11;
wire n_0_58_12;
wire n_0_58_13;
wire n_0_58_14;
wire n_0_58_15;
wire n_0_58_16;
wire n_0_58_17;
wire n_0_58_18;
wire n_0_58_19;
wire n_0_58_20;
wire n_0_58_21;
wire n_0_58_22;
wire n_0_58_23;
wire n_0_58_24;
wire n_0_111;
wire n_0_58_25;
wire n_0_58_26;
wire n_0_58_27;
wire n_0_58_28;
wire n_0_58_29;
wire n_0_58_30;
wire n_0_58_31;
wire n_0_58_32;
wire n_0_58_33;
wire n_0_75_0;
wire n_0_75_1;
wire n_0_75_2;
wire n_0_75_3;
wire n_0_75_4;
wire n_0_75_5;
wire n_0_75_6;
wire n_0_75_7;
wire n_0_75_8;
wire n_0_75_9;
wire n_0_75_10;
wire n_0_75_11;
wire n_0_75_12;
wire n_0_75_13;
wire n_0_75_14;
wire n_0_75_15;
wire n_0_75_16;
wire n_0_75_17;
wire n_0_75_18;
wire n_0_75_19;
wire n_0_75_20;
wire n_0_75_21;
wire n_0_75_22;
wire n_0_75_23;
wire n_0_75_24;
wire n_0_75_25;
wire n_0_75_26;
wire n_0_75_27;
wire n_0_75_28;
wire n_0_75_29;
wire n_0_75_30;
wire n_0_75_31;
wire n_0_75_32;
wire n_0_75_33;
wire n_0_75_34;
wire n_0_112;
wire n_0_113;
wire n_0_92_0;
wire n_0_92_1;
wire n_0_92_2;
wire n_0_92_3;
wire n_0_92_4;
wire n_0_92_5;
wire n_0_92_6;
wire n_0_92_7;
wire n_0_92_8;
wire n_0_92_9;
wire n_0_92_10;
wire n_0_92_11;
wire n_0_92_12;
wire n_0_92_13;
wire n_0_92_14;
wire n_0_92_15;
wire n_0_92_16;
wire n_0_92_17;
wire n_0_92_18;
wire n_0_92_19;
wire n_0_92_20;
wire n_0_92_21;
wire n_0_92_22;
wire n_0_92_23;
wire n_0_92_24;
wire n_0_92_25;
wire n_0_92_26;
wire n_0_114;
wire n_0_109_0;
wire n_0_109_1;
wire n_0_109_2;
wire n_0_109_3;
wire n_0_109_4;
wire n_0_109_5;
wire n_0_109_6;
wire n_0_109_7;
wire n_0_109_8;
wire n_0_109_9;
wire n_0_109_10;
wire n_0_109_11;
wire n_0_109_12;
wire n_0_109_13;
wire n_0_109_14;
wire n_0_109_15;
wire n_0_109_16;
wire n_0_109_17;
wire n_0_109_18;
wire n_0_109_19;
wire n_0_109_20;
wire n_0_109_21;
wire n_0_109_22;
wire n_0_109_23;
wire n_0_109_24;
wire n_0_109_25;
wire n_0_109_26;
wire n_0_109_27;
wire n_0_109_28;
wire n_0_109_29;
wire n_0_109_30;
wire n_0_115;
wire n_0_126_0;
wire n_0_126_1;
wire n_0_126_2;
wire n_0_126_3;
wire n_0_126_4;
wire n_0_126_5;
wire n_0_126_6;
wire n_0_126_7;
wire n_0_126_8;
wire n_0_126_9;
wire n_0_126_10;
wire n_0_126_11;
wire n_0_126_12;
wire n_0_126_13;
wire n_0_126_14;
wire n_0_126_15;
wire n_0_126_16;
wire n_0_126_17;
wire n_0_126_18;
wire n_0_126_19;
wire n_0_126_20;
wire n_0_126_21;
wire n_0_126_22;
wire n_0_126_23;
wire n_0_126_24;
wire n_0_126_25;
wire n_0_126_26;
wire n_0_126_27;
wire n_0_126_28;
wire n_0_126_29;
wire n_0_126_30;
wire n_0_143_0;
wire n_0_143_1;
wire n_0_143_2;
wire n_0_143_3;
wire n_0_143_4;
wire n_0_143_5;
wire n_0_143_6;
wire n_0_143_7;
wire n_0_143_8;
wire n_0_143_9;
wire n_0_143_10;
wire n_0_143_11;
wire n_0_143_12;
wire n_0_143_13;
wire n_0_143_14;
wire n_0_143_15;
wire n_0_143_16;
wire n_0_143_17;
wire n_0_143_18;
wire n_0_143_19;
wire n_0_143_20;
wire n_0_143_21;
wire n_0_143_22;
wire n_0_143_23;
wire n_0_143_24;
wire n_0_143_25;
wire n_0_143_26;
wire n_0_143_27;
wire n_0_143_28;
wire n_0_143_29;
wire n_0_143_30;
wire n_0_143_31;
wire n_0_143_32;
wire n_0_143_33;
wire n_0_143_34;
wire n_0_143_35;
wire n_0_118;
wire n_0_119;
wire n_0_160_0;
wire n_0_160_1;
wire n_0_160_2;
wire n_0_160_3;
wire n_0_160_4;
wire n_0_160_5;
wire n_0_160_6;
wire n_0_160_7;
wire n_0_160_8;
wire n_0_160_9;
wire n_0_160_10;
wire n_0_160_11;
wire n_0_160_12;
wire n_0_160_13;
wire n_0_160_14;
wire n_0_160_15;
wire n_0_160_16;
wire n_0_160_17;
wire n_0_160_18;
wire n_0_160_19;
wire n_0_160_20;
wire n_0_160_21;
wire n_0_160_22;
wire n_0_160_23;
wire n_0_160_24;
wire n_0_160_25;
wire n_0_160_26;
wire n_0_160_27;
wire n_0_160_28;
wire n_0_160_29;
wire n_0_160_30;
wire n_0_177_0;
wire n_0_177_1;
wire n_0_177_2;
wire n_0_177_3;
wire n_0_177_4;
wire n_0_177_5;
wire n_0_177_6;
wire n_0_177_7;
wire n_0_177_8;
wire n_0_177_9;
wire n_0_177_10;
wire n_0_177_11;
wire n_0_177_12;
wire n_0_177_13;
wire n_0_177_14;
wire n_0_177_15;
wire n_0_177_16;
wire n_0_177_17;
wire n_0_177_18;
wire n_0_177_19;
wire n_0_177_20;
wire n_0_177_21;
wire n_0_177_22;
wire n_0_177_23;
wire n_0_177_24;
wire n_0_177_25;
wire n_0_177_26;
wire n_0_177_27;
wire n_0_177_28;
wire n_0_177_29;
wire n_0_177_30;
wire n_0_177_31;
wire n_0_177_32;
wire n_0_177_33;
wire n_0_177_34;
wire n_0_177_35;
wire n_0_120;
wire n_0_135_0;
wire n_0_135_1;
wire n_0_135_2;
wire n_0_135_3;
wire n_0_135_4;
wire n_0_135_5;
wire n_0_135_6;
wire n_0_135_7;
wire n_0_135_8;
wire n_0_135_9;
wire n_0_135_10;
wire n_0_135_11;
wire n_0_135_12;
wire n_0_135_13;
wire n_0_135_14;
wire n_0_135_15;
wire n_0_135_16;
wire n_0_135_17;
wire n_0_135_18;
wire n_0_135_19;
wire n_0_135_20;
wire n_0_135_21;
wire n_0_135_22;
wire n_0_135_23;
wire n_0_135_24;
wire n_0_135_25;
wire n_0_135_26;
wire n_0_135_27;
wire n_0_135_28;
wire n_0_135_29;
wire n_0_135_30;
wire n_0_135_31;
wire n_0_135_32;
wire n_0_135_33;
wire n_0_135_34;
wire n_0_135_35;
wire n_0_121;
wire n_0_2_0;
wire n_0_2_1;
wire n_0_2_2;
wire n_0_2_3;
wire n_0_2_4;
wire n_0_2_5;
wire n_0_2_6;
wire n_0_2_7;
wire n_0_2_8;
wire n_0_2_9;
wire n_0_2_10;
wire n_0_2_11;
wire n_0_2_12;
wire n_0_2_13;
wire n_0_2_14;
wire n_0_2_15;
wire n_0_2_16;
wire n_0_2_17;
wire n_0_2_18;
wire n_0_2_19;
wire n_0_2_20;
wire n_0_2_21;
wire n_0_2_22;
wire n_0_2_23;
wire n_0_2_24;
wire n_0_2_25;
wire n_0_2_26;
wire n_0_2_27;
wire n_0_2_28;
wire n_0_2_29;
wire n_0_2_30;
wire n_0_2_31;
wire n_0_2_32;
wire n_0_2_33;
wire n_0_2_34;
wire n_0_2_35;
wire n_0_2_36;
wire n_0_122;
wire n_0_25_0;
wire n_0_25_1;
wire n_0_25_2;
wire n_0_25_3;
wire n_0_25_4;
wire n_0_25_5;
wire n_0_25_6;
wire n_0_25_7;
wire n_0_25_8;
wire n_0_25_9;
wire n_0_25_10;
wire n_0_25_11;
wire n_0_25_12;
wire n_0_25_13;
wire n_0_25_14;
wire n_0_25_15;
wire n_0_25_16;
wire n_0_25_17;
wire n_0_25_18;
wire n_0_25_19;
wire n_0_25_20;
wire n_0_25_21;
wire n_0_25_22;
wire n_0_25_23;
wire n_0_25_24;
wire n_0_123;
wire n_0_25_25;
wire n_0_25_26;
wire n_0_25_27;
wire n_0_25_28;
wire n_0_25_29;
wire n_0_25_30;
wire n_0_25_31;
wire n_0_25_32;
wire n_0_25_33;
wire n_0_59_0;
wire n_0_59_1;
wire n_0_59_2;
wire n_0_59_3;
wire n_0_59_4;
wire n_0_59_5;
wire n_0_59_6;
wire n_0_59_7;
wire n_0_59_8;
wire n_0_59_9;
wire n_0_59_10;
wire n_0_59_11;
wire n_0_59_12;
wire n_0_59_13;
wire n_0_59_14;
wire n_0_59_15;
wire n_0_59_16;
wire n_0_59_17;
wire n_0_59_18;
wire n_0_59_19;
wire n_0_59_20;
wire n_0_59_21;
wire n_0_59_22;
wire n_0_59_23;
wire n_0_59_24;
wire n_0_124;
wire n_0_59_25;
wire n_0_59_26;
wire n_0_59_27;
wire n_0_59_28;
wire n_0_59_29;
wire n_0_59_30;
wire n_0_59_31;
wire n_0_59_32;
wire n_0_59_33;
wire n_0_76_0;
wire n_0_76_1;
wire n_0_76_2;
wire n_0_76_3;
wire n_0_76_4;
wire n_0_76_5;
wire n_0_76_6;
wire n_0_76_7;
wire n_0_76_8;
wire n_0_76_9;
wire n_0_76_10;
wire n_0_76_11;
wire n_0_76_12;
wire n_0_76_13;
wire n_0_76_14;
wire n_0_76_15;
wire n_0_76_16;
wire n_0_76_17;
wire n_0_76_18;
wire n_0_76_19;
wire n_0_76_20;
wire n_0_76_21;
wire n_0_76_22;
wire n_0_76_23;
wire n_0_76_24;
wire n_0_76_25;
wire n_0_76_26;
wire n_0_76_27;
wire n_0_76_28;
wire n_0_76_29;
wire n_0_76_30;
wire n_0_76_31;
wire n_0_76_32;
wire n_0_76_33;
wire n_0_76_34;
wire n_0_125;
wire n_0_126;
wire n_0_93_0;
wire n_0_93_1;
wire n_0_93_2;
wire n_0_93_3;
wire n_0_93_4;
wire n_0_93_5;
wire n_0_93_6;
wire n_0_93_7;
wire n_0_93_8;
wire n_0_93_9;
wire n_0_93_10;
wire n_0_93_11;
wire n_0_93_12;
wire n_0_93_13;
wire n_0_93_14;
wire n_0_93_15;
wire n_0_93_16;
wire n_0_93_17;
wire n_0_93_18;
wire n_0_93_19;
wire n_0_93_20;
wire n_0_93_21;
wire n_0_93_22;
wire n_0_93_23;
wire n_0_93_24;
wire n_0_93_25;
wire n_0_93_26;
wire n_0_127;
wire n_0_110_0;
wire n_0_110_1;
wire n_0_110_2;
wire n_0_110_3;
wire n_0_110_4;
wire n_0_110_5;
wire n_0_110_6;
wire n_0_110_7;
wire n_0_110_8;
wire n_0_110_9;
wire n_0_110_10;
wire n_0_110_11;
wire n_0_110_12;
wire n_0_110_13;
wire n_0_110_14;
wire n_0_110_15;
wire n_0_110_16;
wire n_0_110_17;
wire n_0_110_18;
wire n_0_110_19;
wire n_0_110_20;
wire n_0_110_21;
wire n_0_110_22;
wire n_0_110_23;
wire n_0_110_24;
wire n_0_110_25;
wire n_0_110_26;
wire n_0_110_27;
wire n_0_110_28;
wire n_0_110_29;
wire n_0_110_30;
wire n_0_128;
wire n_0_127_0;
wire n_0_127_1;
wire n_0_127_2;
wire n_0_127_3;
wire n_0_127_4;
wire n_0_127_5;
wire n_0_127_6;
wire n_0_127_7;
wire n_0_127_8;
wire n_0_127_9;
wire n_0_127_10;
wire n_0_127_11;
wire n_0_127_12;
wire n_0_127_13;
wire n_0_127_14;
wire n_0_127_15;
wire n_0_127_16;
wire n_0_127_17;
wire n_0_127_18;
wire n_0_127_19;
wire n_0_127_20;
wire n_0_127_21;
wire n_0_127_22;
wire n_0_127_23;
wire n_0_127_24;
wire n_0_127_25;
wire n_0_127_26;
wire n_0_127_27;
wire n_0_127_28;
wire n_0_127_29;
wire n_0_127_30;
wire n_0_144_0;
wire n_0_144_1;
wire n_0_144_2;
wire n_0_144_3;
wire n_0_144_4;
wire n_0_144_5;
wire n_0_144_6;
wire n_0_144_7;
wire n_0_144_8;
wire n_0_144_9;
wire n_0_144_10;
wire n_0_144_11;
wire n_0_144_12;
wire n_0_144_13;
wire n_0_144_14;
wire n_0_144_15;
wire n_0_144_16;
wire n_0_144_17;
wire n_0_144_18;
wire n_0_144_19;
wire n_0_144_20;
wire n_0_144_21;
wire n_0_144_22;
wire n_0_144_23;
wire n_0_144_24;
wire n_0_144_25;
wire n_0_144_26;
wire n_0_144_27;
wire n_0_144_28;
wire n_0_144_29;
wire n_0_144_30;
wire n_0_144_31;
wire n_0_144_32;
wire n_0_144_33;
wire n_0_144_34;
wire n_0_144_35;
wire n_0_129;
wire n_0_130;
wire n_0_161_0;
wire n_0_161_1;
wire n_0_161_2;
wire n_0_161_3;
wire n_0_161_4;
wire n_0_161_5;
wire n_0_161_6;
wire n_0_161_7;
wire n_0_161_8;
wire n_0_161_9;
wire n_0_161_10;
wire n_0_161_11;
wire n_0_161_12;
wire n_0_161_13;
wire n_0_161_14;
wire n_0_161_15;
wire n_0_161_16;
wire n_0_161_17;
wire n_0_161_18;
wire n_0_161_19;
wire n_0_161_20;
wire n_0_161_21;
wire n_0_161_22;
wire n_0_161_23;
wire n_0_161_24;
wire n_0_161_25;
wire n_0_161_26;
wire n_0_161_27;
wire n_0_161_28;
wire n_0_161_29;
wire n_0_161_30;
wire n_0_178_0;
wire n_0_178_1;
wire n_0_178_2;
wire n_0_178_3;
wire n_0_178_4;
wire n_0_178_5;
wire n_0_178_6;
wire n_0_178_7;
wire n_0_178_8;
wire n_0_178_9;
wire n_0_178_10;
wire n_0_178_11;
wire n_0_178_12;
wire n_0_178_13;
wire n_0_178_14;
wire n_0_178_15;
wire n_0_178_16;
wire n_0_178_17;
wire n_0_178_18;
wire n_0_178_19;
wire n_0_178_20;
wire n_0_178_21;
wire n_0_178_22;
wire n_0_178_23;
wire n_0_178_24;
wire n_0_178_25;
wire n_0_178_26;
wire n_0_178_27;
wire n_0_178_28;
wire n_0_178_29;
wire n_0_178_30;
wire n_0_178_31;
wire n_0_178_32;
wire n_0_178_33;
wire n_0_178_34;
wire n_0_178_35;
wire n_0_131;
wire n_0_84_0;
wire n_0_84_1;
wire n_0_84_2;
wire n_0_84_3;
wire n_0_84_4;
wire n_0_84_5;
wire n_0_84_6;
wire n_0_84_7;
wire n_0_84_8;
wire n_0_84_9;
wire n_0_84_10;
wire n_0_84_11;
wire n_0_84_12;
wire n_0_84_13;
wire n_0_84_14;
wire n_0_84_15;
wire n_0_84_16;
wire n_0_84_17;
wire n_0_84_18;
wire n_0_84_19;
wire n_0_84_20;
wire n_0_84_21;
wire n_0_84_22;
wire n_0_84_23;
wire n_0_84_24;
wire n_0_84_25;
wire n_0_84_26;
wire n_0_84_27;
wire n_0_84_28;
wire n_0_84_29;
wire n_0_84_30;
wire n_0_84_31;
wire n_0_84_32;
wire n_0_84_33;
wire n_0_84_34;
wire n_0_84_35;
wire n_0_132;
wire n_0_26_0;
wire n_0_26_1;
wire n_0_26_2;
wire n_0_26_3;
wire n_0_26_4;
wire n_0_26_5;
wire n_0_26_6;
wire n_0_26_7;
wire n_0_26_8;
wire n_0_26_9;
wire n_0_26_10;
wire n_0_26_11;
wire n_0_26_12;
wire n_0_26_13;
wire n_0_26_14;
wire n_0_26_15;
wire n_0_26_16;
wire n_0_26_17;
wire n_0_26_18;
wire n_0_26_19;
wire n_0_26_20;
wire n_0_26_21;
wire n_0_26_22;
wire n_0_26_23;
wire n_0_26_24;
wire n_0_26_25;
wire n_0_26_26;
wire n_0_26_27;
wire n_0_26_28;
wire n_0_26_29;
wire n_0_26_30;
wire n_0_26_31;
wire n_0_26_32;
wire n_0_26_33;
wire n_0_26_34;
wire n_0_26_35;
wire n_0_26_36;
wire n_0_133;
wire n_0_43_0;
wire n_0_43_1;
wire n_0_43_2;
wire n_0_43_3;
wire n_0_43_4;
wire n_0_43_5;
wire n_0_43_6;
wire n_0_43_7;
wire n_0_43_8;
wire n_0_43_9;
wire n_0_43_10;
wire n_0_43_11;
wire n_0_43_12;
wire n_0_43_13;
wire n_0_43_14;
wire n_0_43_15;
wire n_0_43_16;
wire n_0_43_17;
wire n_0_43_18;
wire n_0_43_19;
wire n_0_43_20;
wire n_0_43_21;
wire n_0_43_22;
wire n_0_43_23;
wire n_0_43_24;
wire n_0_134;
wire n_0_43_25;
wire n_0_43_26;
wire n_0_43_27;
wire n_0_43_28;
wire n_0_43_29;
wire n_0_43_30;
wire n_0_43_31;
wire n_0_43_32;
wire n_0_43_33;
wire n_0_60_0;
wire n_0_60_1;
wire n_0_60_2;
wire n_0_60_3;
wire n_0_60_4;
wire n_0_60_5;
wire n_0_60_6;
wire n_0_60_7;
wire n_0_60_8;
wire n_0_60_9;
wire n_0_60_10;
wire n_0_60_11;
wire n_0_60_12;
wire n_0_60_13;
wire n_0_60_14;
wire n_0_60_15;
wire n_0_60_16;
wire n_0_60_17;
wire n_0_60_18;
wire n_0_60_19;
wire n_0_60_20;
wire n_0_60_21;
wire n_0_60_22;
wire n_0_60_23;
wire n_0_60_24;
wire n_0_135;
wire n_0_60_25;
wire n_0_60_26;
wire n_0_60_27;
wire n_0_60_28;
wire n_0_60_29;
wire n_0_60_30;
wire n_0_60_31;
wire n_0_60_32;
wire n_0_60_33;
wire n_0_77_0;
wire n_0_77_1;
wire n_0_77_2;
wire n_0_77_3;
wire n_0_77_4;
wire n_0_77_5;
wire n_0_77_6;
wire n_0_77_7;
wire n_0_77_8;
wire n_0_77_9;
wire n_0_77_10;
wire n_0_77_11;
wire n_0_77_12;
wire n_0_77_13;
wire n_0_77_14;
wire n_0_77_15;
wire n_0_77_16;
wire n_0_77_17;
wire n_0_77_18;
wire n_0_77_19;
wire n_0_77_20;
wire n_0_77_21;
wire n_0_77_22;
wire n_0_77_23;
wire n_0_77_24;
wire n_0_77_25;
wire n_0_77_26;
wire n_0_77_27;
wire n_0_77_28;
wire n_0_77_29;
wire n_0_77_30;
wire n_0_77_31;
wire n_0_77_32;
wire n_0_77_33;
wire n_0_77_34;
wire n_0_136;
wire n_0_137;
wire n_0_94_0;
wire n_0_94_1;
wire n_0_94_2;
wire n_0_94_3;
wire n_0_94_4;
wire n_0_94_5;
wire n_0_94_6;
wire n_0_94_7;
wire n_0_94_8;
wire n_0_94_9;
wire n_0_94_10;
wire n_0_94_11;
wire n_0_94_12;
wire n_0_94_13;
wire n_0_94_14;
wire n_0_94_15;
wire n_0_94_16;
wire n_0_94_17;
wire n_0_94_18;
wire n_0_94_19;
wire n_0_94_20;
wire n_0_94_21;
wire n_0_94_22;
wire n_0_94_23;
wire n_0_94_24;
wire n_0_94_25;
wire n_0_94_26;
wire n_0_138;
wire n_0_111_0;
wire n_0_111_1;
wire n_0_111_2;
wire n_0_111_3;
wire n_0_111_4;
wire n_0_111_5;
wire n_0_111_6;
wire n_0_111_7;
wire n_0_111_8;
wire n_0_111_9;
wire n_0_111_10;
wire n_0_111_11;
wire n_0_111_12;
wire n_0_111_13;
wire n_0_111_14;
wire n_0_111_15;
wire n_0_111_16;
wire n_0_111_17;
wire n_0_111_18;
wire n_0_111_19;
wire n_0_111_20;
wire n_0_111_21;
wire n_0_111_22;
wire n_0_111_23;
wire n_0_111_24;
wire n_0_111_25;
wire n_0_111_26;
wire n_0_111_27;
wire n_0_111_28;
wire n_0_111_29;
wire n_0_111_30;
wire n_0_139;
wire n_0_128_0;
wire n_0_128_1;
wire n_0_128_2;
wire n_0_128_3;
wire n_0_128_4;
wire n_0_128_5;
wire n_0_128_6;
wire n_0_128_7;
wire n_0_128_8;
wire n_0_128_9;
wire n_0_128_10;
wire n_0_128_11;
wire n_0_128_12;
wire n_0_128_13;
wire n_0_128_14;
wire n_0_128_15;
wire n_0_128_16;
wire n_0_128_17;
wire n_0_128_18;
wire n_0_128_19;
wire n_0_128_20;
wire n_0_128_21;
wire n_0_128_22;
wire n_0_128_23;
wire n_0_128_24;
wire n_0_128_25;
wire n_0_128_26;
wire n_0_128_27;
wire n_0_128_28;
wire n_0_128_29;
wire n_0_128_30;
wire n_0_145_0;
wire n_0_145_1;
wire n_0_145_2;
wire n_0_145_3;
wire n_0_145_4;
wire n_0_145_5;
wire n_0_145_6;
wire n_0_145_7;
wire n_0_145_8;
wire n_0_145_9;
wire n_0_145_10;
wire n_0_145_11;
wire n_0_145_12;
wire n_0_145_13;
wire n_0_145_14;
wire n_0_145_15;
wire n_0_145_16;
wire n_0_145_17;
wire n_0_145_18;
wire n_0_145_19;
wire n_0_145_20;
wire n_0_145_21;
wire n_0_145_22;
wire n_0_145_23;
wire n_0_145_24;
wire n_0_145_25;
wire n_0_145_26;
wire n_0_145_27;
wire n_0_145_28;
wire n_0_145_29;
wire n_0_145_30;
wire n_0_145_31;
wire n_0_145_32;
wire n_0_145_33;
wire n_0_145_34;
wire n_0_145_35;
wire n_0_140;
wire n_0_141;
wire n_0_162_0;
wire n_0_162_1;
wire n_0_162_2;
wire n_0_162_3;
wire n_0_162_4;
wire n_0_162_5;
wire n_0_162_6;
wire n_0_162_7;
wire n_0_162_8;
wire n_0_162_9;
wire n_0_162_10;
wire n_0_162_11;
wire n_0_162_12;
wire n_0_162_13;
wire n_0_162_14;
wire n_0_162_15;
wire n_0_162_16;
wire n_0_162_17;
wire n_0_162_18;
wire n_0_162_19;
wire n_0_162_20;
wire n_0_162_21;
wire n_0_162_22;
wire n_0_162_23;
wire n_0_162_24;
wire n_0_162_25;
wire n_0_162_26;
wire n_0_162_27;
wire n_0_162_28;
wire n_0_162_29;
wire n_0_162_30;
wire n_0_179_0;
wire n_0_179_1;
wire n_0_179_2;
wire n_0_179_3;
wire n_0_179_4;
wire n_0_179_5;
wire n_0_179_6;
wire n_0_179_7;
wire n_0_179_8;
wire n_0_179_9;
wire n_0_179_10;
wire n_0_179_11;
wire n_0_179_12;
wire n_0_179_13;
wire n_0_179_14;
wire n_0_179_15;
wire n_0_179_16;
wire n_0_179_17;
wire n_0_179_18;
wire n_0_179_19;
wire n_0_179_20;
wire n_0_179_21;
wire n_0_179_22;
wire n_0_179_23;
wire n_0_179_24;
wire n_0_179_25;
wire n_0_179_26;
wire n_0_179_27;
wire n_0_179_28;
wire n_0_179_29;
wire n_0_179_30;
wire n_0_179_31;
wire n_0_179_32;
wire n_0_179_33;
wire n_0_179_34;
wire n_0_179_35;
wire n_0_142;
wire n_0_42_0;
wire n_0_42_1;
wire n_0_42_2;
wire n_0_42_3;
wire n_0_42_4;
wire n_0_42_5;
wire n_0_42_6;
wire n_0_42_7;
wire n_0_42_8;
wire n_0_42_9;
wire n_0_42_10;
wire n_0_42_11;
wire n_0_42_12;
wire n_0_42_13;
wire n_0_42_14;
wire n_0_42_15;
wire n_0_42_16;
wire n_0_42_17;
wire n_0_42_18;
wire n_0_42_19;
wire n_0_42_20;
wire n_0_42_21;
wire n_0_42_22;
wire n_0_42_23;
wire n_0_42_24;
wire n_0_42_25;
wire n_0_42_26;
wire n_0_42_27;
wire n_0_42_28;
wire n_0_42_29;
wire n_0_42_30;
wire n_0_42_31;
wire n_0_42_32;
wire n_0_42_33;
wire n_0_42_34;
wire n_0_42_35;
wire n_0_143;
wire n_0_27_0;
wire n_0_27_1;
wire n_0_27_2;
wire n_0_27_3;
wire n_0_27_4;
wire n_0_27_5;
wire n_0_27_6;
wire n_0_27_7;
wire n_0_27_8;
wire n_0_27_9;
wire n_0_27_10;
wire n_0_27_11;
wire n_0_27_12;
wire n_0_27_13;
wire n_0_27_14;
wire n_0_27_15;
wire n_0_27_16;
wire n_0_27_17;
wire n_0_27_18;
wire n_0_27_19;
wire n_0_27_20;
wire n_0_27_21;
wire n_0_27_22;
wire n_0_27_23;
wire n_0_27_24;
wire n_0_27_25;
wire n_0_27_26;
wire n_0_27_27;
wire n_0_27_28;
wire n_0_27_29;
wire n_0_27_30;
wire n_0_27_31;
wire n_0_27_32;
wire n_0_27_33;
wire n_0_27_34;
wire n_0_27_35;
wire n_0_27_36;
wire n_0_144;
wire n_0_44_0;
wire n_0_44_1;
wire n_0_44_2;
wire n_0_44_3;
wire n_0_44_4;
wire n_0_44_5;
wire n_0_44_6;
wire n_0_44_7;
wire n_0_44_8;
wire n_0_44_9;
wire n_0_44_10;
wire n_0_44_11;
wire n_0_44_12;
wire n_0_44_13;
wire n_0_44_14;
wire n_0_44_15;
wire n_0_44_16;
wire n_0_44_17;
wire n_0_44_18;
wire n_0_44_19;
wire n_0_44_20;
wire n_0_44_21;
wire n_0_44_22;
wire n_0_44_23;
wire n_0_44_24;
wire n_0_145;
wire n_0_44_25;
wire n_0_44_26;
wire n_0_44_27;
wire n_0_44_28;
wire n_0_44_29;
wire n_0_44_30;
wire n_0_44_31;
wire n_0_44_32;
wire n_0_44_33;
wire n_0_61_0;
wire n_0_61_1;
wire n_0_61_2;
wire n_0_61_3;
wire n_0_61_4;
wire n_0_61_5;
wire n_0_61_6;
wire n_0_61_7;
wire n_0_61_8;
wire n_0_61_9;
wire n_0_61_10;
wire n_0_61_11;
wire n_0_61_12;
wire n_0_61_13;
wire n_0_61_14;
wire n_0_61_15;
wire n_0_61_16;
wire n_0_61_17;
wire n_0_61_18;
wire n_0_61_19;
wire n_0_61_20;
wire n_0_61_21;
wire n_0_61_22;
wire n_0_61_23;
wire n_0_61_24;
wire n_0_146;
wire n_0_61_25;
wire n_0_61_26;
wire n_0_61_27;
wire n_0_61_28;
wire n_0_61_29;
wire n_0_61_30;
wire n_0_61_31;
wire n_0_61_32;
wire n_0_61_33;
wire n_0_78_0;
wire n_0_78_1;
wire n_0_78_2;
wire n_0_78_3;
wire n_0_78_4;
wire n_0_78_5;
wire n_0_78_6;
wire n_0_78_7;
wire n_0_78_8;
wire n_0_78_9;
wire n_0_78_10;
wire n_0_78_11;
wire n_0_78_12;
wire n_0_78_13;
wire n_0_78_14;
wire n_0_78_15;
wire n_0_78_16;
wire n_0_78_17;
wire n_0_78_18;
wire n_0_78_19;
wire n_0_78_20;
wire n_0_78_21;
wire n_0_78_22;
wire n_0_78_23;
wire n_0_78_24;
wire n_0_78_25;
wire n_0_78_26;
wire n_0_78_27;
wire n_0_78_28;
wire n_0_78_29;
wire n_0_78_30;
wire n_0_78_31;
wire n_0_78_32;
wire n_0_78_33;
wire n_0_78_34;
wire n_0_147;
wire n_0_148;
wire n_0_95_0;
wire n_0_95_1;
wire n_0_95_2;
wire n_0_95_3;
wire n_0_95_4;
wire n_0_95_5;
wire n_0_95_6;
wire n_0_95_7;
wire n_0_95_8;
wire n_0_95_9;
wire n_0_95_10;
wire n_0_95_11;
wire n_0_95_12;
wire n_0_95_13;
wire n_0_95_14;
wire n_0_95_15;
wire n_0_95_16;
wire n_0_95_17;
wire n_0_95_18;
wire n_0_95_19;
wire n_0_95_20;
wire n_0_95_21;
wire n_0_95_22;
wire n_0_95_23;
wire n_0_95_24;
wire n_0_95_25;
wire n_0_95_26;
wire n_0_149;
wire n_0_112_0;
wire n_0_112_1;
wire n_0_112_2;
wire n_0_112_3;
wire n_0_112_4;
wire n_0_112_5;
wire n_0_112_6;
wire n_0_112_7;
wire n_0_112_8;
wire n_0_112_9;
wire n_0_112_10;
wire n_0_112_11;
wire n_0_112_12;
wire n_0_112_13;
wire n_0_112_14;
wire n_0_112_15;
wire n_0_112_16;
wire n_0_112_17;
wire n_0_112_18;
wire n_0_112_19;
wire n_0_112_20;
wire n_0_112_21;
wire n_0_112_22;
wire n_0_112_23;
wire n_0_112_24;
wire n_0_112_25;
wire n_0_112_26;
wire n_0_112_27;
wire n_0_112_28;
wire n_0_112_29;
wire n_0_112_30;
wire n_0_152;
wire n_0_129_0;
wire n_0_129_1;
wire n_0_129_2;
wire n_0_129_3;
wire n_0_129_4;
wire n_0_129_5;
wire n_0_129_6;
wire n_0_129_7;
wire n_0_129_8;
wire n_0_129_9;
wire n_0_129_10;
wire n_0_129_11;
wire n_0_129_12;
wire n_0_129_13;
wire n_0_129_14;
wire n_0_129_15;
wire n_0_129_16;
wire n_0_129_17;
wire n_0_129_18;
wire n_0_129_19;
wire n_0_129_20;
wire n_0_129_21;
wire n_0_129_22;
wire n_0_129_23;
wire n_0_129_24;
wire n_0_129_25;
wire n_0_129_26;
wire n_0_129_27;
wire n_0_129_28;
wire n_0_129_29;
wire n_0_129_30;
wire n_0_146_0;
wire n_0_146_1;
wire n_0_146_2;
wire n_0_146_3;
wire n_0_146_4;
wire n_0_146_5;
wire n_0_146_6;
wire n_0_146_7;
wire n_0_146_8;
wire n_0_146_9;
wire n_0_146_10;
wire n_0_146_11;
wire n_0_146_12;
wire n_0_146_13;
wire n_0_146_14;
wire n_0_146_15;
wire n_0_146_16;
wire n_0_146_17;
wire n_0_146_18;
wire n_0_146_19;
wire n_0_146_20;
wire n_0_146_21;
wire n_0_146_22;
wire n_0_146_23;
wire n_0_146_24;
wire n_0_146_25;
wire n_0_146_26;
wire n_0_146_27;
wire n_0_146_28;
wire n_0_146_29;
wire n_0_146_30;
wire n_0_146_31;
wire n_0_146_32;
wire n_0_146_33;
wire n_0_146_34;
wire n_0_146_35;
wire n_0_153;
wire n_0_154;
wire n_0_163_0;
wire n_0_163_1;
wire n_0_163_2;
wire n_0_163_3;
wire n_0_163_4;
wire n_0_163_5;
wire n_0_163_6;
wire n_0_163_7;
wire n_0_163_8;
wire n_0_163_9;
wire n_0_163_10;
wire n_0_163_11;
wire n_0_163_12;
wire n_0_163_13;
wire n_0_163_14;
wire n_0_163_15;
wire n_0_163_16;
wire n_0_163_17;
wire n_0_163_18;
wire n_0_163_19;
wire n_0_163_20;
wire n_0_163_21;
wire n_0_163_22;
wire n_0_163_23;
wire n_0_163_24;
wire n_0_163_25;
wire n_0_163_26;
wire n_0_163_27;
wire n_0_163_28;
wire n_0_163_29;
wire n_0_163_30;
wire n_0_180_0;
wire n_0_180_1;
wire n_0_180_2;
wire n_0_180_3;
wire n_0_180_4;
wire n_0_180_5;
wire n_0_180_6;
wire n_0_180_7;
wire n_0_180_8;
wire n_0_180_9;
wire n_0_180_10;
wire n_0_180_11;
wire n_0_180_12;
wire n_0_180_13;
wire n_0_180_14;
wire n_0_180_15;
wire n_0_180_16;
wire n_0_180_17;
wire n_0_180_18;
wire n_0_180_19;
wire n_0_180_20;
wire n_0_180_21;
wire n_0_180_22;
wire n_0_180_23;
wire n_0_180_24;
wire n_0_180_25;
wire n_0_180_26;
wire n_0_180_27;
wire n_0_180_28;
wire n_0_180_29;
wire n_0_180_30;
wire n_0_180_31;
wire n_0_180_32;
wire n_0_180_33;
wire n_0_180_34;
wire n_0_180_35;
wire n_0_155;
wire n_0_152_0;
wire n_0_152_1;
wire n_0_152_2;
wire n_0_152_3;
wire n_0_152_4;
wire n_0_152_5;
wire n_0_152_6;
wire n_0_152_7;
wire n_0_152_8;
wire n_0_152_9;
wire n_0_152_10;
wire n_0_152_11;
wire n_0_152_12;
wire n_0_152_13;
wire n_0_152_14;
wire n_0_152_15;
wire n_0_152_16;
wire n_0_152_17;
wire n_0_152_18;
wire n_0_152_19;
wire n_0_152_20;
wire n_0_152_21;
wire n_0_152_22;
wire n_0_152_23;
wire n_0_152_24;
wire n_0_152_25;
wire n_0_152_26;
wire n_0_152_27;
wire n_0_152_28;
wire n_0_152_29;
wire n_0_152_30;
wire n_0_152_31;
wire n_0_152_32;
wire n_0_152_33;
wire n_0_152_34;
wire n_0_152_35;
wire n_0_156;
wire n_0_28_0;
wire n_0_28_1;
wire n_0_28_2;
wire n_0_28_3;
wire n_0_28_4;
wire n_0_28_5;
wire n_0_28_6;
wire n_0_28_7;
wire n_0_28_8;
wire n_0_28_9;
wire n_0_28_10;
wire n_0_28_11;
wire n_0_28_12;
wire n_0_28_13;
wire n_0_28_14;
wire n_0_28_15;
wire n_0_28_16;
wire n_0_28_17;
wire n_0_28_18;
wire n_0_28_19;
wire n_0_28_20;
wire n_0_28_21;
wire n_0_28_22;
wire n_0_28_23;
wire n_0_28_24;
wire n_0_28_25;
wire n_0_28_26;
wire n_0_28_27;
wire n_0_28_28;
wire n_0_28_29;
wire n_0_28_30;
wire n_0_28_31;
wire n_0_28_32;
wire n_0_28_33;
wire n_0_28_34;
wire n_0_28_35;
wire n_0_28_36;
wire n_0_157;
wire n_0_45_0;
wire n_0_45_1;
wire n_0_45_2;
wire n_0_45_3;
wire n_0_45_4;
wire n_0_45_5;
wire n_0_45_6;
wire n_0_45_7;
wire n_0_45_8;
wire n_0_45_9;
wire n_0_45_10;
wire n_0_45_11;
wire n_0_45_12;
wire n_0_45_13;
wire n_0_45_14;
wire n_0_45_15;
wire n_0_45_16;
wire n_0_45_17;
wire n_0_45_18;
wire n_0_45_19;
wire n_0_45_20;
wire n_0_45_21;
wire n_0_45_22;
wire n_0_45_23;
wire n_0_45_24;
wire n_0_158;
wire n_0_45_25;
wire n_0_45_26;
wire n_0_45_27;
wire n_0_45_28;
wire n_0_45_29;
wire n_0_45_30;
wire n_0_45_31;
wire n_0_45_32;
wire n_0_45_33;
wire n_0_62_0;
wire n_0_62_1;
wire n_0_62_2;
wire n_0_62_3;
wire n_0_62_4;
wire n_0_62_5;
wire n_0_62_6;
wire n_0_62_7;
wire n_0_62_8;
wire n_0_62_9;
wire n_0_62_10;
wire n_0_62_11;
wire n_0_62_12;
wire n_0_62_13;
wire n_0_62_14;
wire n_0_62_15;
wire n_0_62_16;
wire n_0_62_17;
wire n_0_62_18;
wire n_0_62_19;
wire n_0_62_20;
wire n_0_62_21;
wire n_0_62_22;
wire n_0_62_23;
wire n_0_62_24;
wire n_0_159;
wire n_0_62_25;
wire n_0_62_26;
wire n_0_62_27;
wire n_0_62_28;
wire n_0_62_29;
wire n_0_62_30;
wire n_0_62_31;
wire n_0_62_32;
wire n_0_62_33;
wire n_0_63_0;
wire n_0_63_1;
wire n_0_63_2;
wire n_0_63_3;
wire n_0_63_4;
wire n_0_63_5;
wire n_0_63_6;
wire n_0_63_7;
wire n_0_63_8;
wire n_0_63_9;
wire n_0_63_10;
wire n_0_63_11;
wire n_0_63_12;
wire n_0_63_13;
wire n_0_63_14;
wire n_0_63_15;
wire n_0_63_16;
wire n_0_63_17;
wire n_0_63_18;
wire n_0_63_19;
wire n_0_63_20;
wire n_0_63_21;
wire n_0_63_22;
wire n_0_63_23;
wire n_0_63_24;
wire n_0_63_25;
wire n_0_63_26;
wire n_0_63_27;
wire n_0_63_28;
wire n_0_63_29;
wire n_0_63_30;
wire n_0_63_31;
wire n_0_63_32;
wire n_0_63_33;
wire n_0_63_34;
wire n_0_160;
wire n_0_79_0;
wire n_0_79_1;
wire n_0_79_2;
wire n_0_79_3;
wire n_0_79_4;
wire n_0_79_5;
wire n_0_79_6;
wire n_0_79_7;
wire n_0_79_8;
wire n_0_79_9;
wire n_0_79_10;
wire n_0_79_11;
wire n_0_79_12;
wire n_0_79_13;
wire n_0_79_14;
wire n_0_79_15;
wire n_0_79_16;
wire n_0_79_17;
wire n_0_79_18;
wire n_0_79_19;
wire n_0_79_20;
wire n_0_79_21;
wire n_0_79_22;
wire n_0_79_23;
wire n_0_79_24;
wire n_0_79_25;
wire n_0_79_26;
wire n_0_79_27;
wire n_0_79_28;
wire n_0_79_29;
wire n_0_79_30;
wire n_0_79_31;
wire n_0_79_32;
wire n_0_79_33;
wire n_0_79_34;
wire n_0_161;
wire n_0_162;
wire n_0_80_0;
wire n_0_80_1;
wire n_0_80_2;
wire n_0_80_3;
wire n_0_80_4;
wire n_0_80_5;
wire n_0_80_6;
wire n_0_80_7;
wire n_0_80_8;
wire n_0_80_9;
wire n_0_80_10;
wire n_0_80_11;
wire n_0_80_12;
wire n_0_80_13;
wire n_0_80_14;
wire n_0_80_15;
wire n_0_80_16;
wire n_0_80_17;
wire n_0_80_18;
wire n_0_80_19;
wire n_0_80_20;
wire n_0_80_21;
wire n_0_80_22;
wire n_0_80_23;
wire n_0_80_24;
wire n_0_80_25;
wire n_0_80_26;
wire n_0_163;
wire n_0_81_0;
wire n_0_81_1;
wire n_0_81_2;
wire n_0_81_3;
wire n_0_81_4;
wire n_0_81_5;
wire n_0_81_6;
wire n_0_81_7;
wire n_0_81_8;
wire n_0_81_9;
wire n_0_81_10;
wire n_0_81_11;
wire n_0_81_12;
wire n_0_81_13;
wire n_0_81_14;
wire n_0_81_15;
wire n_0_81_16;
wire n_0_81_17;
wire n_0_81_18;
wire n_0_81_19;
wire n_0_81_20;
wire n_0_81_21;
wire n_0_81_22;
wire n_0_81_23;
wire n_0_81_24;
wire n_0_81_25;
wire n_0_81_26;
wire n_0_164;
wire n_0_96_0;
wire n_0_96_1;
wire n_0_96_2;
wire n_0_96_3;
wire n_0_96_4;
wire n_0_96_5;
wire n_0_96_6;
wire n_0_96_7;
wire n_0_96_8;
wire n_0_96_9;
wire n_0_96_10;
wire n_0_96_11;
wire n_0_96_12;
wire n_0_96_13;
wire n_0_96_14;
wire n_0_96_15;
wire n_0_96_16;
wire n_0_96_17;
wire n_0_96_18;
wire n_0_96_19;
wire n_0_96_20;
wire n_0_96_21;
wire n_0_96_22;
wire n_0_96_23;
wire n_0_96_24;
wire n_0_96_25;
wire n_0_96_26;
wire n_0_165;
wire n_0_113_0;
wire n_0_113_1;
wire n_0_113_2;
wire n_0_113_3;
wire n_0_113_4;
wire n_0_113_5;
wire n_0_113_6;
wire n_0_113_7;
wire n_0_113_8;
wire n_0_113_9;
wire n_0_113_10;
wire n_0_113_11;
wire n_0_113_12;
wire n_0_113_13;
wire n_0_113_14;
wire n_0_113_15;
wire n_0_113_16;
wire n_0_113_17;
wire n_0_113_18;
wire n_0_113_19;
wire n_0_113_20;
wire n_0_113_21;
wire n_0_113_22;
wire n_0_113_23;
wire n_0_113_24;
wire n_0_113_25;
wire n_0_113_26;
wire n_0_113_27;
wire n_0_113_28;
wire n_0_113_29;
wire n_0_113_30;
wire n_0_166;
wire n_0_130_0;
wire n_0_130_1;
wire n_0_130_2;
wire n_0_130_3;
wire n_0_130_4;
wire n_0_130_5;
wire n_0_130_6;
wire n_0_130_7;
wire n_0_130_8;
wire n_0_130_9;
wire n_0_130_10;
wire n_0_130_11;
wire n_0_130_12;
wire n_0_130_13;
wire n_0_130_14;
wire n_0_130_15;
wire n_0_130_16;
wire n_0_130_17;
wire n_0_130_18;
wire n_0_130_19;
wire n_0_130_20;
wire n_0_130_21;
wire n_0_130_22;
wire n_0_130_23;
wire n_0_130_24;
wire n_0_130_25;
wire n_0_130_26;
wire n_0_130_27;
wire n_0_130_28;
wire n_0_130_29;
wire n_0_130_30;
wire n_0_131_0;
wire n_0_131_1;
wire n_0_131_2;
wire n_0_131_3;
wire n_0_131_4;
wire n_0_131_5;
wire n_0_131_6;
wire n_0_131_7;
wire n_0_131_8;
wire n_0_131_9;
wire n_0_131_10;
wire n_0_131_11;
wire n_0_131_12;
wire n_0_131_13;
wire n_0_131_14;
wire n_0_131_15;
wire n_0_131_16;
wire n_0_131_17;
wire n_0_131_18;
wire n_0_131_19;
wire n_0_131_20;
wire n_0_131_21;
wire n_0_131_22;
wire n_0_131_23;
wire n_0_131_24;
wire n_0_131_25;
wire n_0_131_26;
wire n_0_131_27;
wire n_0_131_28;
wire n_0_131_29;
wire n_0_131_30;
wire n_0_131_31;
wire n_0_131_32;
wire n_0_131_33;
wire n_0_131_34;
wire n_0_131_35;
wire n_0_167;
wire n_0_132_0;
wire n_0_132_1;
wire n_0_132_2;
wire n_0_132_3;
wire n_0_132_4;
wire n_0_132_5;
wire n_0_132_6;
wire n_0_132_7;
wire n_0_132_8;
wire n_0_132_9;
wire n_0_132_10;
wire n_0_132_11;
wire n_0_132_12;
wire n_0_132_13;
wire n_0_132_14;
wire n_0_132_15;
wire n_0_132_16;
wire n_0_132_17;
wire n_0_132_18;
wire n_0_132_19;
wire n_0_132_20;
wire n_0_132_21;
wire n_0_132_22;
wire n_0_132_23;
wire n_0_132_24;
wire n_0_132_25;
wire n_0_132_26;
wire n_0_132_27;
wire n_0_132_28;
wire n_0_132_29;
wire n_0_132_30;
wire n_0_132_31;
wire n_0_132_32;
wire n_0_132_33;
wire n_0_132_34;
wire n_0_132_35;
wire n_0_168;
wire n_0_147_0;
wire n_0_147_1;
wire n_0_147_2;
wire n_0_147_3;
wire n_0_147_4;
wire n_0_147_5;
wire n_0_147_6;
wire n_0_147_7;
wire n_0_147_8;
wire n_0_147_9;
wire n_0_147_10;
wire n_0_147_11;
wire n_0_147_12;
wire n_0_147_13;
wire n_0_147_14;
wire n_0_147_15;
wire n_0_147_16;
wire n_0_147_17;
wire n_0_147_18;
wire n_0_147_19;
wire n_0_147_20;
wire n_0_147_21;
wire n_0_147_22;
wire n_0_147_23;
wire n_0_147_24;
wire n_0_147_25;
wire n_0_147_26;
wire n_0_147_27;
wire n_0_147_28;
wire n_0_147_29;
wire n_0_147_30;
wire n_0_147_31;
wire n_0_147_32;
wire n_0_147_33;
wire n_0_147_34;
wire n_0_147_35;
wire n_0_169;
wire n_0_170;
wire n_0_164_0;
wire n_0_164_1;
wire n_0_164_2;
wire n_0_164_3;
wire n_0_164_4;
wire n_0_164_5;
wire n_0_164_6;
wire n_0_164_7;
wire n_0_164_8;
wire n_0_164_9;
wire n_0_164_10;
wire n_0_164_11;
wire n_0_164_12;
wire n_0_164_13;
wire n_0_164_14;
wire n_0_164_15;
wire n_0_164_16;
wire n_0_164_17;
wire n_0_164_18;
wire n_0_164_19;
wire n_0_164_20;
wire n_0_164_21;
wire n_0_164_22;
wire n_0_164_23;
wire n_0_164_24;
wire n_0_164_25;
wire n_0_164_26;
wire n_0_164_27;
wire n_0_164_28;
wire n_0_164_29;
wire n_0_164_30;
wire n_0_165_0;
wire n_0_165_1;
wire n_0_165_2;
wire n_0_165_3;
wire n_0_165_4;
wire n_0_165_5;
wire n_0_165_6;
wire n_0_165_7;
wire n_0_165_8;
wire n_0_165_9;
wire n_0_165_10;
wire n_0_165_11;
wire n_0_165_12;
wire n_0_165_13;
wire n_0_165_14;
wire n_0_165_15;
wire n_0_165_16;
wire n_0_165_17;
wire n_0_165_18;
wire n_0_165_19;
wire n_0_165_20;
wire n_0_165_21;
wire n_0_165_22;
wire n_0_165_23;
wire n_0_165_24;
wire n_0_165_25;
wire n_0_165_26;
wire n_0_165_27;
wire n_0_165_28;
wire n_0_165_29;
wire n_0_165_30;
wire n_0_165_31;
wire n_0_165_32;
wire n_0_165_33;
wire n_0_165_34;
wire n_0_165_35;
wire n_0_171;
wire n_0_166_0;
wire n_0_166_1;
wire n_0_166_2;
wire n_0_166_3;
wire n_0_166_4;
wire n_0_166_5;
wire n_0_166_6;
wire n_0_166_7;
wire n_0_166_8;
wire n_0_166_9;
wire n_0_166_10;
wire n_0_166_11;
wire n_0_166_12;
wire n_0_166_13;
wire n_0_166_14;
wire n_0_166_15;
wire n_0_166_16;
wire n_0_166_17;
wire n_0_166_18;
wire n_0_166_19;
wire n_0_166_20;
wire n_0_166_21;
wire n_0_166_22;
wire n_0_166_23;
wire n_0_166_24;
wire n_0_166_25;
wire n_0_166_26;
wire n_0_166_27;
wire n_0_166_28;
wire n_0_166_29;
wire n_0_166_30;
wire n_0_166_31;
wire n_0_166_32;
wire n_0_166_33;
wire n_0_166_34;
wire n_0_166_35;
wire n_0_172;
wire n_0_181_0;
wire n_0_181_1;
wire n_0_181_2;
wire n_0_181_3;
wire n_0_181_4;
wire n_0_181_5;
wire n_0_181_6;
wire n_0_181_7;
wire n_0_181_8;
wire n_0_181_9;
wire n_0_181_10;
wire n_0_181_11;
wire n_0_181_12;
wire n_0_181_13;
wire n_0_181_14;
wire n_0_181_15;
wire n_0_181_16;
wire n_0_181_17;
wire n_0_181_18;
wire n_0_181_19;
wire n_0_181_20;
wire n_0_181_21;
wire n_0_181_22;
wire n_0_181_23;
wire n_0_181_24;
wire n_0_181_25;
wire n_0_181_26;
wire n_0_181_27;
wire n_0_181_28;
wire n_0_181_29;
wire n_0_181_30;
wire n_0_181_31;
wire n_0_181_32;
wire n_0_181_33;
wire n_0_181_34;
wire n_0_181_35;
wire n_0_173;
wire n_0_182_0;
wire n_0_182_1;
wire n_0_182_2;
wire n_0_182_3;
wire n_0_182_4;
wire n_0_182_5;
wire n_0_182_6;
wire n_0_182_7;
wire n_0_182_8;
wire n_0_182_9;
wire n_0_182_10;
wire n_0_182_11;
wire n_0_182_12;
wire n_0_182_13;
wire n_0_182_14;
wire n_0_182_15;
wire n_0_182_16;
wire n_0_182_17;
wire n_0_182_18;
wire n_0_182_19;
wire n_0_182_20;
wire n_0_182_21;
wire n_0_182_22;
wire n_0_182_23;
wire n_0_182_24;
wire n_0_182_25;
wire n_0_182_26;
wire n_0_182_27;
wire n_0_182_28;
wire n_0_182_29;
wire n_0_182_30;
wire n_0_182_31;
wire n_0_182_32;
wire n_0_182_33;
wire n_0_182_34;
wire n_0_182_35;
wire n_0_174;
wire n_0_183_0;
wire n_0_183_1;
wire n_0_183_2;
wire n_0_183_3;
wire n_0_183_4;
wire n_0_183_5;
wire n_0_183_6;
wire n_0_183_7;
wire n_0_183_8;
wire n_0_183_9;
wire n_0_183_10;
wire n_0_183_11;
wire n_0_183_12;
wire n_0_183_13;
wire n_0_183_14;
wire n_0_183_15;
wire n_0_183_16;
wire n_0_183_17;
wire n_0_183_18;
wire n_0_183_19;
wire n_0_183_20;
wire n_0_183_21;
wire n_0_183_22;
wire n_0_183_23;
wire n_0_183_24;
wire n_0_183_25;
wire n_0_183_26;
wire n_0_183_27;
wire n_0_183_28;
wire n_0_183_29;
wire n_0_183_30;
wire n_0_183_31;
wire n_0_183_32;
wire n_0_183_33;
wire n_0_183_34;
wire n_0_183_35;
wire n_0_175;
wire n_0_169_0;
wire n_0_169_1;
wire n_0_169_2;
wire n_0_169_3;
wire n_0_169_4;
wire n_0_169_5;
wire n_0_169_6;
wire n_0_169_7;
wire n_0_169_8;
wire n_0_169_9;
wire n_0_169_10;
wire n_0_169_11;
wire n_0_169_12;
wire n_0_169_13;
wire n_0_169_14;
wire n_0_169_15;
wire n_0_169_16;
wire n_0_169_17;
wire n_0_169_18;
wire n_0_169_19;
wire n_0_169_20;
wire n_0_169_21;
wire n_0_169_22;
wire n_0_169_23;
wire n_0_169_24;
wire n_0_169_25;
wire n_0_169_26;
wire n_0_169_27;
wire n_0_169_28;
wire n_0_169_29;
wire n_0_169_30;
wire n_0_169_31;
wire n_0_169_32;
wire n_0_169_33;
wire n_0_169_34;
wire n_0_169_35;
wire n_0_176;
wire n_0_197_0;
wire n_0_197_1;
wire n_0_197_2;
wire n_0_197_3;
wire n_0_197_4;
wire n_0_197_5;
wire n_0_197_6;
wire n_0_197_7;
wire n_0_197_8;
wire n_0_197_9;
wire n_0_197_10;
wire n_0_197_11;
wire n_0_197_12;
wire n_0_197_13;
wire n_0_197_14;
wire n_0_197_15;
wire n_0_197_16;
wire n_0_197_17;
wire n_0_197_18;
wire n_0_197_19;
wire n_0_197_20;
wire n_0_197_21;
wire n_0_197_22;
wire n_0_197_23;
wire n_0_197_24;
wire n_0_197_25;
wire n_0_197_26;
wire n_0_197_27;
wire n_0_197_28;
wire n_0_197_29;
wire n_0_197_30;
wire n_0_197_31;
wire n_0_197_32;
wire n_0_197_33;
wire n_0_197_34;
wire n_0_197_35;
wire n_0_197_36;
wire n_0_177;
wire n_0_198_0;
wire n_0_198_1;
wire n_0_198_2;
wire n_0_198_3;
wire n_0_198_4;
wire n_0_198_5;
wire n_0_198_6;
wire n_0_198_7;
wire n_0_198_8;
wire n_0_198_9;
wire n_0_198_10;
wire n_0_198_11;
wire n_0_198_12;
wire n_0_198_13;
wire n_0_198_14;
wire n_0_198_15;
wire n_0_198_16;
wire n_0_198_17;
wire n_0_198_18;
wire n_0_198_19;
wire n_0_198_20;
wire n_0_198_21;
wire n_0_198_22;
wire n_0_198_23;
wire n_0_198_24;
wire n_0_198_25;
wire n_0_198_26;
wire n_0_198_27;
wire n_0_198_28;
wire n_0_198_29;
wire n_0_198_30;
wire n_0_198_31;
wire n_0_198_32;
wire n_0_198_33;
wire n_0_198_34;
wire n_0_198_35;
wire n_0_198_36;
wire n_0_178;
wire n_0_64_0;
wire n_0_64_1;
wire n_0_64_2;
wire n_0_64_3;
wire n_0_64_4;
wire n_0_64_5;
wire n_0_64_6;
wire n_0_64_7;
wire n_0_64_8;
wire n_0_64_9;
wire n_0_64_10;
wire n_0_64_11;
wire n_0_64_12;
wire n_0_64_13;
wire n_0_64_14;
wire n_0_64_15;
wire n_0_64_16;
wire n_0_64_17;
wire n_0_64_18;
wire n_0_64_19;
wire n_0_64_20;
wire n_0_64_21;
wire n_0_64_22;
wire n_0_64_23;
wire n_0_64_24;
wire n_0_64_25;
wire n_0_64_26;
wire n_0_64_27;
wire n_0_64_28;
wire n_0_64_29;
wire n_0_64_30;
wire n_0_64_31;
wire n_0_64_32;
wire n_0_64_33;
wire n_0_64_34;
wire n_0_64_35;
wire n_0_64_36;
wire n_0_179;
wire n_0_133_0;
wire n_0_133_1;
wire n_0_133_2;
wire n_0_133_3;
wire n_0_133_4;
wire n_0_133_5;
wire n_0_133_6;
wire n_0_133_7;
wire n_0_133_8;
wire n_0_133_9;
wire n_0_133_10;
wire n_0_133_11;
wire n_0_133_12;
wire n_0_133_13;
wire n_0_133_14;
wire n_0_133_15;
wire n_0_133_16;
wire n_0_133_17;
wire n_0_133_18;
wire n_0_133_19;
wire n_0_133_20;
wire n_0_133_21;
wire n_0_133_22;
wire n_0_133_23;
wire n_0_133_24;
wire n_0_133_25;
wire n_0_133_26;
wire n_0_133_27;
wire n_0_133_28;
wire n_0_133_29;
wire n_0_133_30;
wire n_0_133_31;
wire n_0_133_32;
wire n_0_133_33;
wire n_0_133_34;
wire n_0_180;
wire n_0_167_0;
wire n_0_167_1;
wire n_0_167_2;
wire n_0_167_3;
wire n_0_167_4;
wire n_0_167_5;
wire n_0_167_6;
wire n_0_167_7;
wire n_0_167_8;
wire n_0_167_9;
wire n_0_167_10;
wire n_0_167_11;
wire n_0_167_12;
wire n_0_167_13;
wire n_0_167_14;
wire n_0_167_15;
wire n_0_167_16;
wire n_0_167_17;
wire n_0_167_18;
wire n_0_167_19;
wire n_0_167_20;
wire n_0_167_21;
wire n_0_167_22;
wire n_0_167_23;
wire n_0_167_24;
wire n_0_167_25;
wire n_0_167_26;
wire n_0_167_27;
wire n_0_167_28;
wire n_0_167_29;
wire n_0_167_30;
wire n_0_167_31;
wire n_0_167_32;
wire n_0_167_33;
wire n_0_167_34;
wire n_0_167_35;
wire n_0_181;
wire n_0_184_0;
wire n_0_184_1;
wire n_0_184_2;
wire n_0_184_3;
wire n_0_184_4;
wire n_0_184_5;
wire n_0_184_6;
wire n_0_184_7;
wire n_0_184_8;
wire n_0_184_9;
wire n_0_184_10;
wire n_0_184_11;
wire n_0_184_12;
wire n_0_184_13;
wire n_0_184_14;
wire n_0_184_15;
wire n_0_184_16;
wire n_0_184_17;
wire n_0_184_18;
wire n_0_184_19;
wire n_0_184_20;
wire n_0_184_21;
wire n_0_184_22;
wire n_0_184_23;
wire n_0_184_24;
wire n_0_184_25;
wire n_0_184_26;
wire n_0_184_27;
wire n_0_184_28;
wire n_0_184_29;
wire n_0_184_30;
wire n_0_184_31;
wire n_0_184_32;
wire n_0_184_33;
wire n_0_184_34;
wire n_0_184_35;
wire n_0_182;
wire n_0_188_0;
wire n_0_188_1;
wire n_0_188_2;
wire n_0_188_3;
wire n_0_188_4;
wire n_0_188_5;
wire n_0_188_6;
wire n_0_188_7;
wire n_0_188_8;
wire n_0_188_9;
wire n_0_188_10;
wire n_0_188_11;
wire n_0_188_12;
wire n_0_188_13;
wire n_0_188_14;
wire n_0_188_15;
wire n_0_188_16;
wire n_0_188_17;
wire n_0_188_18;
wire n_0_188_19;
wire n_0_188_20;
wire n_0_188_21;
wire n_0_188_22;
wire n_0_188_23;
wire n_0_188_24;
wire n_0_188_25;
wire n_0_188_26;
wire n_0_188_27;
wire n_0_188_28;
wire n_0_188_29;
wire n_0_188_30;
wire n_0_188_31;
wire n_0_188_32;
wire n_0_188_33;
wire n_0_188_34;
wire n_0_188_35;
wire n_0_183;
wire n_0_65_0;
wire n_0_65_1;
wire n_0_65_2;
wire n_0_65_3;
wire n_0_65_4;
wire n_0_65_5;
wire n_0_65_6;
wire n_0_65_7;
wire n_0_65_8;
wire n_0_65_9;
wire n_0_65_10;
wire n_0_65_11;
wire n_0_65_12;
wire n_0_65_13;
wire n_0_65_14;
wire n_0_65_15;
wire n_0_65_16;
wire n_0_65_17;
wire n_0_65_18;
wire n_0_65_19;
wire n_0_65_20;
wire n_0_65_21;
wire n_0_65_22;
wire n_0_65_23;
wire n_0_65_24;
wire n_0_65_25;
wire n_0_65_26;
wire n_0_65_27;
wire n_0_65_28;
wire n_0_65_29;
wire n_0_65_30;
wire n_0_65_31;
wire n_0_65_32;
wire n_0_65_33;
wire n_0_65_34;
wire n_0_65_35;
wire n_0_65_36;
wire n_0_184;
wire n_0_82_0;
wire n_0_82_1;
wire n_0_82_2;
wire n_0_82_3;
wire n_0_82_4;
wire n_0_82_5;
wire n_0_82_6;
wire n_0_82_7;
wire n_0_82_8;
wire n_0_82_9;
wire n_0_82_10;
wire n_0_82_11;
wire n_0_82_12;
wire n_0_82_13;
wire n_0_82_14;
wire n_0_82_15;
wire n_0_82_16;
wire n_0_82_17;
wire n_0_82_18;
wire n_0_82_19;
wire n_0_82_20;
wire n_0_82_21;
wire n_0_82_22;
wire n_0_82_23;
wire n_0_82_24;
wire n_0_82_25;
wire n_0_82_26;
wire n_0_82_27;
wire n_0_82_28;
wire n_0_82_29;
wire n_0_82_30;
wire n_0_82_31;
wire n_0_82_32;
wire n_0_82_33;
wire n_0_82_34;
wire n_0_186;
wire n_0_188;
wire n_0_29_0;
wire n_0_29_1;
wire n_0_29_2;
wire n_0_29_3;
wire n_0_29_4;
wire n_0_29_5;
wire n_0_29_6;
wire n_0_29_7;
wire n_0_29_8;
wire n_0_29_9;
wire n_0_29_10;
wire n_0_29_11;
wire n_0_29_12;
wire n_0_29_13;
wire n_0_29_14;
wire n_0_29_15;
wire n_0_29_16;
wire n_0_29_17;
wire n_0_29_18;
wire n_0_29_19;
wire n_0_29_20;
wire n_0_29_21;
wire n_0_29_22;
wire n_0_29_23;
wire n_0_29_24;
wire n_0_29_25;
wire n_0_29_26;
wire n_0_46_0;
wire n_0_46_1;
wire n_0_46_2;
wire n_0_46_3;
wire n_0_46_4;
wire n_0_46_5;
wire n_0_46_6;
wire n_0_46_7;
wire n_0_46_8;
wire n_0_46_9;
wire n_0_46_10;
wire n_0_46_11;
wire n_0_46_12;
wire n_0_46_13;
wire n_0_46_14;
wire n_0_46_15;
wire n_0_46_16;
wire n_0_46_17;
wire n_0_46_18;
wire n_0_46_19;
wire n_0_46_20;
wire n_0_46_21;
wire n_0_46_22;
wire n_0_46_23;
wire n_0_46_24;
wire n_0_189;
wire n_0_46_25;
wire n_0_46_26;
wire n_0_46_27;
wire n_0_46_28;
wire n_0_46_29;
wire n_0_46_30;
wire n_0_46_31;
wire n_0_46_32;
wire n_0_46_33;
wire n_0_97_0;
wire n_0_97_1;
wire n_0_97_2;
wire n_0_97_3;
wire n_0_97_4;
wire n_0_97_5;
wire n_0_97_6;
wire n_0_97_7;
wire n_0_97_8;
wire n_0_97_9;
wire n_0_97_10;
wire n_0_97_11;
wire n_0_97_12;
wire n_0_97_13;
wire n_0_97_14;
wire n_0_97_15;
wire n_0_97_16;
wire n_0_97_17;
wire n_0_97_18;
wire n_0_97_19;
wire n_0_97_20;
wire n_0_97_21;
wire n_0_97_22;
wire n_0_97_23;
wire n_0_97_24;
wire n_0_190;
wire n_0_97_25;
wire n_0_97_26;
wire n_0_97_27;
wire n_0_97_28;
wire n_0_97_29;
wire n_0_97_30;
wire n_0_97_31;
wire n_0_97_32;
wire n_0_97_33;
wire n_0_191;
wire n_0_114_0;
wire n_0_114_1;
wire n_0_114_2;
wire n_0_114_3;
wire n_0_114_4;
wire n_0_114_5;
wire n_0_114_6;
wire n_0_114_7;
wire n_0_114_8;
wire n_0_114_9;
wire n_0_114_10;
wire n_0_114_11;
wire n_0_114_12;
wire n_0_114_13;
wire n_0_114_14;
wire n_0_114_15;
wire n_0_114_16;
wire n_0_114_17;
wire n_0_114_18;
wire n_0_114_19;
wire n_0_114_20;
wire n_0_114_21;
wire n_0_114_22;
wire n_0_114_23;
wire n_0_114_24;
wire n_0_114_25;
wire n_0_114_26;
wire n_0_114_27;
wire n_0_114_28;
wire n_0_114_29;
wire n_0_114_30;
wire n_0_192;
wire n_0_148_0;
wire n_0_148_1;
wire n_0_148_2;
wire n_0_148_3;
wire n_0_148_4;
wire n_0_148_5;
wire n_0_148_6;
wire n_0_148_7;
wire n_0_148_8;
wire n_0_148_9;
wire n_0_148_10;
wire n_0_148_11;
wire n_0_148_12;
wire n_0_148_13;
wire n_0_148_14;
wire n_0_148_15;
wire n_0_148_16;
wire n_0_148_17;
wire n_0_148_18;
wire n_0_148_19;
wire n_0_148_20;
wire n_0_148_21;
wire n_0_148_22;
wire n_0_148_23;
wire n_0_148_24;
wire n_0_148_25;
wire n_0_148_26;
wire n_0_148_27;
wire n_0_148_28;
wire n_0_148_29;
wire n_0_148_30;
wire n_0_193;
wire n_0_83_0;
wire n_0_83_1;
wire n_0_83_2;
wire n_0_83_3;
wire n_0_83_4;
wire n_0_83_5;
wire n_0_83_6;
wire n_0_83_7;
wire n_0_83_8;
wire n_0_83_9;
wire n_0_83_10;
wire n_0_83_11;
wire n_0_83_12;
wire n_0_83_13;
wire n_0_83_14;
wire n_0_83_15;
wire n_0_83_16;
wire n_0_83_17;
wire n_0_83_18;
wire n_0_83_19;
wire n_0_83_20;
wire n_0_83_21;
wire n_0_83_22;
wire n_0_83_23;
wire n_0_83_24;
wire n_0_83_25;
wire n_0_83_26;
wire n_0_83_27;
wire n_0_83_28;
wire n_0_83_29;
wire n_0_83_30;
wire n_0_194;
wire n_0_186_0;
wire n_0_186_6;
wire n_0_186_7;
wire n_0_186_8;
wire n_0_186_9;
wire n_0_186_10;
wire n_0_186_11;
wire n_0_186_12;
wire n_0_186_27;
wire n_0_186_28;
wire n_0_186_1;
wire n_0_186_2;
wire n_0_186_13;
wire n_0_186_3;
wire n_0_186_4;
wire n_0_186_5;
wire n_0_186_14;
wire n_0_186_15;
wire n_0_186_16;
wire n_0_186_17;
wire n_0_186_18;
wire n_0_186_19;
wire n_0_186_20;
wire n_0_186_21;
wire n_0_186_22;
wire n_0_186_23;
wire n_0_186_24;
wire n_0_186_25;
wire n_0_186_26;
wire n_0_168_0;
wire n_0_168_1;
wire n_0_168_2;
wire n_0_168_3;
wire n_0_168_4;
wire n_0_168_5;
wire n_0_168_6;
wire n_0_168_7;
wire n_0_168_8;
wire n_0_168_9;
wire n_0_168_10;
wire n_0_168_11;
wire n_0_168_12;
wire n_0_168_13;
wire n_0_168_14;
wire n_0_168_15;
wire n_0_168_16;
wire n_0_168_17;
wire n_0_168_18;
wire n_0_168_19;
wire n_0_168_20;
wire n_0_168_21;
wire n_0_168_22;
wire n_0_168_23;
wire n_0_168_24;
wire n_0_168_25;
wire n_0_168_26;
wire n_0_168_27;
wire n_0_168_28;
wire n_0_168_29;
wire n_0_168_30;
wire n_0_168_31;
wire n_0_168_32;
wire n_0_168_33;
wire n_0_168_34;
wire n_0_168_35;
wire n_0_195;
wire n_0_185_0;
wire n_0_185_1;
wire n_0_185_2;
wire n_0_185_3;
wire n_0_185_4;
wire n_0_185_5;
wire n_0_185_6;
wire n_0_185_7;
wire n_0_185_8;
wire n_0_185_9;
wire n_0_185_10;
wire n_0_185_11;
wire n_0_185_12;
wire n_0_185_13;
wire n_0_185_14;
wire n_0_185_15;
wire n_0_185_16;
wire n_0_185_17;
wire n_0_185_18;
wire n_0_185_19;
wire n_0_185_20;
wire n_0_185_21;
wire n_0_185_22;
wire n_0_185_23;
wire n_0_185_24;
wire n_0_185_25;
wire n_0_185_26;
wire n_0_185_27;
wire n_0_185_28;
wire n_0_185_29;
wire n_0_185_30;
wire n_0_185_31;
wire n_0_185_32;
wire n_0_185_33;
wire n_0_185_34;
wire n_0_185_35;
wire n_0_196;
wire n_0_30_0;
wire n_0_30_1;
wire n_0_30_2;
wire n_0_30_3;
wire n_0_30_4;
wire n_0_30_5;
wire n_0_30_6;
wire n_0_30_7;
wire n_0_30_8;
wire n_0_30_9;
wire n_0_30_10;
wire n_0_30_11;
wire n_0_30_12;
wire n_0_30_13;
wire n_0_30_14;
wire n_0_30_15;
wire n_0_30_16;
wire n_0_30_17;
wire n_0_30_18;
wire n_0_30_19;
wire n_0_30_20;
wire n_0_30_21;
wire n_0_30_22;
wire n_0_30_23;
wire n_0_30_24;
wire n_0_30_25;
wire n_0_30_26;
wire n_0_30_27;
wire n_0_30_28;
wire n_0_30_29;
wire n_0_30_30;
wire n_0_30_31;
wire n_0_30_32;
wire n_0_30_33;
wire n_0_30_34;
wire n_0_30_35;
wire n_0_197;
wire n_0_47_0;
wire n_0_47_1;
wire n_0_47_2;
wire n_0_47_3;
wire n_0_47_4;
wire n_0_47_5;
wire n_0_47_6;
wire n_0_47_7;
wire n_0_47_8;
wire n_0_47_9;
wire n_0_47_10;
wire n_0_47_11;
wire n_0_47_12;
wire n_0_47_13;
wire n_0_47_14;
wire n_0_47_15;
wire n_0_47_16;
wire n_0_47_17;
wire n_0_47_18;
wire n_0_47_19;
wire n_0_47_20;
wire n_0_47_21;
wire n_0_47_22;
wire n_0_47_23;
wire n_0_47_24;
wire n_0_198;
wire n_0_47_25;
wire n_0_47_26;
wire n_0_47_27;
wire n_0_47_28;
wire n_0_47_29;
wire n_0_47_30;
wire n_0_47_31;
wire n_0_47_32;
wire n_0_47_33;
wire n_0_98_0;
wire n_0_98_1;
wire n_0_98_2;
wire n_0_98_3;
wire n_0_98_4;
wire n_0_98_5;
wire n_0_98_6;
wire n_0_98_7;
wire n_0_98_8;
wire n_0_98_9;
wire n_0_98_10;
wire n_0_98_11;
wire n_0_98_12;
wire n_0_98_13;
wire n_0_98_14;
wire n_0_98_15;
wire n_0_98_16;
wire n_0_98_17;
wire n_0_98_18;
wire n_0_98_19;
wire n_0_98_20;
wire n_0_98_21;
wire n_0_98_22;
wire n_0_98_23;
wire n_0_98_24;
wire n_0_0;
wire n_0_98_25;
wire n_0_98_26;
wire n_0_98_27;
wire n_0_98_28;
wire n_0_98_29;
wire n_0_98_30;
wire n_0_98_31;
wire n_0_98_32;
wire n_0_98_33;
wire n_0_1;
wire n_0_115_0;
wire n_0_115_1;
wire n_0_115_2;
wire n_0_115_3;
wire n_0_115_4;
wire n_0_115_5;
wire n_0_115_6;
wire n_0_115_7;
wire n_0_115_8;
wire n_0_115_9;
wire n_0_115_10;
wire n_0_115_11;
wire n_0_115_12;
wire n_0_115_13;
wire n_0_115_14;
wire n_0_115_15;
wire n_0_115_16;
wire n_0_115_17;
wire n_0_115_18;
wire n_0_115_19;
wire n_0_115_20;
wire n_0_115_21;
wire n_0_115_22;
wire n_0_115_23;
wire n_0_115_24;
wire n_0_115_25;
wire n_0_115_26;
wire n_0_115_27;
wire n_0_115_28;
wire n_0_115_29;
wire n_0_115_30;
wire n_0_2;
wire n_0_134_0;
wire n_0_134_1;
wire n_0_134_2;
wire n_0_134_3;
wire n_0_134_4;
wire n_0_134_5;
wire n_0_134_6;
wire n_0_134_7;
wire n_0_134_8;
wire n_0_134_9;
wire n_0_134_10;
wire n_0_134_11;
wire n_0_134_12;
wire n_0_134_13;
wire n_0_134_14;
wire n_0_134_15;
wire n_0_134_16;
wire n_0_134_17;
wire n_0_134_18;
wire n_0_134_19;
wire n_0_134_20;
wire n_0_134_21;
wire n_0_134_22;
wire n_0_134_23;
wire n_0_134_24;
wire n_0_134_25;
wire n_0_134_26;
wire n_0_134_27;
wire n_0_134_28;
wire n_0_134_29;
wire n_0_134_30;
wire n_0_3;
wire n_0_193_0;
wire n_0_193_1;
wire n_0_193_2;
wire n_0_193_3;
wire n_0_193_4;
wire n_0_193_5;
wire n_0_193_6;
wire n_0_193_7;
wire n_0_193_8;
wire n_0_193_9;
wire n_0_193_10;
wire n_0_193_11;
wire n_0_193_12;
wire n_0_193_13;
wire n_0_193_14;
wire n_0_193_15;
wire n_0_193_16;
wire n_0_193_17;
wire n_0_193_18;
wire n_0_193_19;
wire n_0_193_20;
wire n_0_193_21;
wire n_0_193_22;
wire n_0_193_23;
wire n_0_193_24;
wire n_0_193_25;
wire n_0_193_26;
wire n_0_193_27;
wire n_0_193_28;
wire n_0_193_29;
wire n_0_193_30;
wire n_0_49;
wire n_0_99_0;
wire n_0_99_1;
wire n_0_99_2;
wire n_0_99_3;
wire n_0_99_4;
wire n_0_99_5;
wire n_0_99_6;
wire n_0_99_7;
wire n_0_99_8;
wire n_0_99_9;
wire n_0_99_10;
wire n_0_99_11;
wire n_0_99_12;
wire n_0_99_13;
wire n_0_99_14;
wire n_0_99_15;
wire n_0_99_16;
wire n_0_99_17;
wire n_0_99_18;
wire n_0_99_19;
wire n_0_99_20;
wire n_0_99_21;
wire n_0_99_22;
wire n_0_99_23;
wire n_0_99_24;
wire n_0_99_25;
wire n_0_99_26;
wire n_0_99_27;
wire n_0_99_28;
wire n_0_99_29;
wire n_0_99_30;
wire n_0_116_0;
wire n_0_116_1;
wire n_0_116_2;
wire n_0_116_3;
wire n_0_116_4;
wire n_0_116_5;
wire n_0_116_6;
wire n_0_116_7;
wire n_0_116_8;
wire n_0_116_9;
wire n_0_116_10;
wire n_0_116_11;
wire n_0_116_12;
wire n_0_116_13;
wire n_0_116_14;
wire n_0_116_15;
wire n_0_116_16;
wire n_0_116_17;
wire n_0_116_18;
wire n_0_116_19;
wire n_0_116_20;
wire n_0_116_21;
wire n_0_116_22;
wire n_0_116_23;
wire n_0_116_24;
wire n_0_116_25;
wire n_0_116_26;
wire n_0_116_27;
wire n_0_116_28;
wire n_0_116_29;
wire n_0_116_30;
wire n_0_65;
wire n_0_66;
wire n_0_149_0;
wire n_0_149_1;
wire n_0_149_2;
wire n_0_149_3;
wire n_0_149_4;
wire n_0_149_5;
wire n_0_149_6;
wire n_0_149_7;
wire n_0_149_8;
wire n_0_149_9;
wire n_0_149_10;
wire n_0_149_11;
wire n_0_149_12;
wire n_0_149_13;
wire n_0_149_14;
wire n_0_149_15;
wire n_0_149_16;
wire n_0_149_17;
wire n_0_149_18;
wire n_0_149_19;
wire n_0_149_20;
wire n_0_149_21;
wire n_0_149_22;
wire n_0_149_23;
wire n_0_149_24;
wire n_0_149_25;
wire n_0_149_26;
wire n_0_149_27;
wire n_0_149_28;
wire n_0_149_29;
wire n_0_149_30;
wire n_0_150_0;
wire n_0_150_1;
wire n_0_150_2;
wire n_0_150_3;
wire n_0_150_4;
wire n_0_150_5;
wire n_0_150_6;
wire n_0_150_7;
wire n_0_150_8;
wire n_0_150_9;
wire n_0_150_10;
wire n_0_150_11;
wire n_0_150_12;
wire n_0_150_13;
wire n_0_150_14;
wire n_0_150_15;
wire n_0_150_16;
wire n_0_150_17;
wire n_0_150_18;
wire n_0_150_19;
wire n_0_150_20;
wire n_0_150_21;
wire n_0_150_22;
wire n_0_150_23;
wire n_0_150_24;
wire n_0_150_25;
wire n_0_150_26;
wire n_0_150_27;
wire n_0_150_28;
wire n_0_150_29;
wire n_0_150_30;
wire n_0_99;
wire n_0_100;
wire n_0_31_0;
wire n_0_31_1;
wire n_0_31_2;
wire n_0_31_3;
wire n_0_31_4;
wire n_0_31_5;
wire n_0_31_6;
wire n_0_31_7;
wire n_0_31_8;
wire n_0_31_9;
wire n_0_31_10;
wire n_0_31_11;
wire n_0_31_12;
wire n_0_31_13;
wire n_0_31_14;
wire n_0_31_15;
wire n_0_31_16;
wire n_0_31_17;
wire n_0_31_18;
wire n_0_31_19;
wire n_0_31_20;
wire n_0_31_21;
wire n_0_31_22;
wire n_0_31_23;
wire n_0_31_24;
wire n_0_31_25;
wire n_0_31_26;
wire n_0_31_27;
wire n_0_31_28;
wire n_0_31_29;
wire n_0_31_30;
wire n_0_187_0;
wire n_0_187_1;
wire n_0_187_2;
wire n_0_187_3;
wire n_0_187_4;
wire n_0_187_5;
wire n_0_187_6;
wire n_0_187_7;
wire n_0_187_8;
wire n_0_187_9;
wire n_0_187_10;
wire n_0_187_11;
wire n_0_187_12;
wire n_0_187_13;
wire n_0_187_14;
wire n_0_187_15;
wire n_0_187_16;
wire n_0_187_17;
wire n_0_187_18;
wire n_0_187_19;
wire n_0_187_20;
wire n_0_187_21;
wire n_0_187_22;
wire n_0_187_23;
wire n_0_187_24;
wire n_0_187_25;
wire n_0_187_26;
wire n_0_187_27;
wire n_0_187_28;
wire n_0_187_29;
wire n_0_187_30;
wire n_0_116;
wire n_0_48_0;
wire n_0_48_1;
wire n_0_48_2;
wire n_0_48_3;
wire n_0_48_4;
wire n_0_48_5;
wire n_0_48_6;
wire n_0_48_7;
wire n_0_48_8;
wire n_0_48_9;
wire n_0_48_10;
wire n_0_48_11;
wire n_0_48_12;
wire n_0_48_13;
wire n_0_48_14;
wire n_0_48_15;
wire n_0_48_16;
wire n_0_48_17;
wire n_0_48_18;
wire n_0_48_19;
wire n_0_48_20;
wire n_0_48_21;
wire n_0_48_22;
wire n_0_48_23;
wire n_0_48_24;
wire n_0_117;
wire n_0_48_25;
wire n_0_48_26;
wire n_0_48_27;
wire n_0_48_28;
wire n_0_48_29;
wire n_0_48_30;
wire n_0_48_31;
wire n_0_48_32;
wire n_0_48_33;
wire n_0_6_0;
wire n_0_6_1;
wire n_0_6_2;
wire n_0_6_3;
wire n_0_6_4;
wire n_0_6_5;
wire n_0_6_6;
wire n_0_6_7;
wire n_0_6_8;
wire n_0_6_9;
wire n_0_6_10;
wire n_0_6_11;
wire n_0_6_12;
wire n_0_6_13;
wire n_0_6_14;
wire n_0_6_15;
wire n_0_6_16;
wire n_0_6_17;
wire n_0_6_18;
wire n_0_6_19;
wire n_0_6_20;
wire n_0_6_21;
wire n_0_6_22;
wire n_0_6_23;
wire n_0_6_24;
wire n_0_150;
wire n_0_6_25;
wire n_0_6_26;
wire n_0_6_27;
wire n_0_6_28;
wire n_0_6_29;
wire n_0_6_30;
wire n_0_6_31;
wire n_0_6_32;
wire n_0_6_33;
wire n_0_190_0;
wire n_0_190_1;
wire n_0_190_2;
wire n_0_190_3;
wire n_0_190_4;
wire n_0_190_5;
wire n_0_151;
wire n_0_190_6;
wire n_0_190_7;
wire n_0_190_8;
wire n_0_190_9;
wire n_0_190_10;
wire n_0_190_11;
wire n_0_190_12;
wire n_0_190_13;
wire n_0_190_14;
wire n_0_190_15;
wire n_0_190_16;
wire n_0_190_17;
wire n_0_190_18;
wire n_0_190_19;
wire n_0_190_20;
wire n_0_190_21;
wire n_0_190_22;
wire n_0_190_23;
wire n_0_190_24;
wire n_0_190_25;
wire n_0_190_26;
wire n_0_190_27;
wire n_0_190_28;
wire n_0_190_29;
wire n_0_190_30;
wire n_0_190_31;
wire n_0_190_32;
wire n_0_190_33;
wire n_0_190_34;
wire n_0_190_35;
wire n_0_190_36;
wire n_0_190_37;
wire n_0_190_38;
wire n_0_32_0;
wire n_0_32_1;
wire n_0_32_2;
wire n_0_32_3;
wire n_0_32_4;
wire n_0_32_5;
wire n_0_32_6;
wire n_0_32_7;
wire n_0_32_8;
wire n_0_32_9;
wire n_0_32_10;
wire n_0_32_11;
wire n_0_32_12;
wire n_0_32_13;
wire n_0_32_14;
wire n_0_32_15;
wire n_0_32_16;
wire n_0_32_17;
wire n_0_32_18;
wire n_0_32_19;
wire n_0_32_20;
wire n_0_32_21;
wire n_0_32_22;
wire n_0_32_23;
wire n_0_32_24;
wire n_0_185;
wire n_0_32_25;
wire n_0_32_26;
wire n_0_32_27;
wire n_0_32_28;
wire n_0_32_29;
wire n_0_32_30;
wire n_0_32_31;
wire n_0_32_32;
wire n_0_32_33;
wire n_0_7_0;
wire n_0_7_1;
wire n_0_7_2;
wire n_0_7_3;
wire n_0_7_4;
wire n_0_7_5;
wire n_0_7_6;
wire n_0_7_7;
wire n_0_7_8;
wire n_0_7_9;
wire n_0_187;
wire n_0_7_10;
wire n_0_7_11;
wire n_0_7_12;
wire n_0_7_13;
wire n_0_7_14;
wire n_0_7_15;
wire n_0_7_16;
wire n_0_7_17;
wire n_0_7_18;
wire n_0_7_19;
wire n_0_7_20;
wire n_0_7_21;
wire n_0_7_22;
wire n_0_7_23;
wire n_0_7_24;
wire n_0_7_25;
wire n_0_7_26;
wire n_0_7_27;
wire n_0_7_28;
wire n_0_7_29;
wire n_0_7_30;
wire n_0_7_31;
wire n_0_7_32;
wire n_0_7_33;
wire n_0_7_34;
wire n_0_7_35;
wire n_0_7_36;
wire n_0_7_37;
wire n_0_7_38;
wire n_0_49_0;
wire n_0_49_1;
wire n_0_49_2;
wire n_0_49_3;
wire n_0_49_4;
wire n_0_49_5;
wire n_0_4;
wire n_0_49_6;
wire n_0_49_7;
wire n_0_49_8;
wire n_0_49_9;
wire n_0_49_10;
wire n_0_49_11;
wire n_0_49_12;
wire n_0_49_13;
wire n_0_49_14;
wire n_0_49_15;
wire n_0_49_16;
wire n_0_49_17;
wire n_0_49_18;
wire n_0_49_19;
wire n_0_49_20;
wire n_0_49_21;
wire n_0_49_22;
wire n_0_49_23;
wire n_0_49_24;
wire n_0_49_25;
wire n_0_49_26;
wire n_0_49_27;
wire n_0_49_28;
wire n_0_49_29;
wire n_0_49_30;
wire n_0_49_31;
wire n_0_49_32;
wire n_0_49_33;
wire n_0_49_34;
wire n_0_49_35;
wire n_0_49_36;
wire n_0_49_37;
wire n_0_49_38;
wire n_0_5;
wire n_0_66_0;
wire n_0_66_1;
wire n_0_189_0;
wire n_0_189_1;
wire n_0_189_2;
wire n_0_189_3;
wire n_0_189_4;
wire n_0_189_5;
wire n_0_189_6;
wire n_0_189_7;
wire n_0_189_8;
wire n_0_189_9;
wire n_0_189_10;
wire n_0_189_11;
wire n_0_189_12;
wire n_0_189_13;
wire n_0_189_14;
wire n_0_189_15;
wire n_0_189_16;
wire n_0_189_17;
wire n_0_189_18;
wire n_0_189_19;
wire n_0_189_20;
wire n_0_189_21;
wire n_0_189_22;
wire n_0_189_23;
wire n_0_189_24;
wire n_0_189_25;
wire n_0_189_26;
wire n_0_189_27;
wire n_0_189_28;
wire n_0_6;
wire n_0_189_29;
wire n_0_189_30;
wire n_0_189_31;
wire n_0_189_32;
wire n_0_189_33;
wire n_0_189_34;
wire n_0_189_35;
wire n_0_1_0;
wire n_0_1_1;
wire n_0_1_2;
wire n_0_1_3;
wire n_0_1_4;
wire n_0_1_5;
wire n_0_1_6;
wire n_0_1_7;
wire n_0_1_8;
wire n_0_1_9;
wire n_0_1_10;
wire n_0_1_11;
wire n_0_1_12;
wire n_0_1_13;
wire n_0_1_14;
wire n_0_1_15;
wire n_0_1_16;
wire n_0_1_17;
wire n_0_1_18;
wire n_0_1_19;
wire n_0_1_20;
wire n_0_1_21;
wire n_0_1_22;
wire n_0_1_23;
wire n_0_1_24;
wire n_0_1_25;
wire n_0_1_26;
wire n_0_1_27;
wire n_0_1_28;
wire n_0_1_29;
wire n_0_1_30;
wire n_0_1_31;
wire n_0_1_32;
wire n_0_1_33;
wire n_0_1_34;
wire n_0_1_35;
wire n_0_1_36;
wire n_0_7;
wire n_0_72;
wire n_0_4_0;
wire n_0_4_1;
wire n_0_11;
wire n_0_4_2;
wire n_0_4_3;
wire n_0_73;
wire n_0_4_4;
wire n_0_4_5;
wire n_0_9;
wire n_0_4_6;
wire n_0_4_7;
wire n_0_74;
wire n_0_4_8;
wire n_0_4_9;
wire n_0_8;
wire n_0_4_10;
wire n_0_4_11;
wire n_0_4_12;
wire n_0_4_13;
wire n_0_4_14;
wire n_0_4_15;
wire n_0_4_16;
wire n_0_4_17;
wire n_0_4_18;
wire n_0_4_19;
wire n_0_4_20;
wire n_0_4_21;
wire n_0_4_22;
wire n_0_4_23;
wire n_0_4_24;
wire n_0_4_25;
wire n_0_4_26;
wire n_0_4_27;
wire n_0_4_28;
wire n_0_4_29;
wire n_0_4_30;
wire n_0_4_31;
wire n_0_4_32;
wire n_0_4_33;
wire n_0_4_34;
wire n_0_4_35;
wire n_0_4_36;
wire n_0_4_37;
wire n_0_4_38;
wire n_0_4_39;
wire n_0_4_40;
wire n_0_4_41;
wire n_0_4_42;
wire n_0_4_43;
wire n_0_4_44;
wire n_0_4_45;
wire n_0_4_46;
wire n_0_4_47;
wire n_0_4_48;
wire n_0_4_49;
wire n_0_4_50;
wire n_0_4_51;
wire n_0_4_52;
wire n_0_4_53;
wire n_0_4_54;
wire n_0_4_55;
wire n_0_4_56;
wire n_0_4_57;
wire n_0_4_58;
wire n_0_4_59;
wire n_0_4_60;
wire n_0_4_61;
wire n_0_4_62;
wire n_0_4_63;
wire n_0_4_64;
wire n_0_4_65;
wire n_0_4_89;
wire n_0_4_66;
wire n_0_4_67;
wire n_0_4_68;
wire n_0_4_93;
wire n_0_4_69;
wire n_0_4_70;
wire n_0_4_71;
wire n_0_4_72;
wire n_0_4_73;
wire n_0_4_74;
wire n_0_4_75;
wire n_0_4_76;
wire n_0_4_77;
wire n_0_4_78;
wire n_0_4_79;
wire n_0_4_105;
wire n_0_4_80;
wire n_0_4_81;
wire n_0_4_82;
wire n_0_4_109;
wire n_0_4_83;
wire n_0_4_84;
wire n_0_4_85;
wire n_0_4_86;
wire n_0_4_87;
wire n_0_4_88;
wire n_0_4_253;
wire n_0_4_90;
wire n_0_4_91;
wire n_0_4_92;
wire n_0_4_254;
wire n_0_4_94;
wire n_0_4_95;
wire n_0_4_96;
wire n_0_4_97;
wire n_0_4_98;
wire n_0_4_99;
wire n_0_4_100;
wire n_0_4_101;
wire n_0_4_102;
wire n_0_4_103;
wire n_0_4_104;
wire n_0_4_255;
wire n_0_4_106;
wire n_0_4_107;
wire n_0_4_108;
wire n_0_4_256;
wire n_0_4_110;
wire n_0_4_111;
wire n_0_4_112;
wire n_0_4_113;
wire n_0_4_114;
wire n_0_4_115;
wire n_0_4_139;
wire n_0_4_116;
wire n_0_4_117;
wire n_0_4_118;
wire n_0_4_140;
wire n_0_4_119;
wire n_0_4_120;
wire n_0_4_121;
wire n_0_4_122;
wire n_0_4_123;
wire n_0_4_124;
wire n_0_4_125;
wire n_0_4_126;
wire n_0_4_127;
wire n_0_4_128;
wire n_0_4_129;
wire n_0_4_144;
wire n_0_4_130;
wire n_0_4_131;
wire n_0_4_132;
wire n_0_4_156;
wire n_0_4_133;
wire n_0_4_134;
wire n_0_4_135;
wire n_0_4_136;
wire n_0_4_137;
wire n_0_4_138;
wire n_0_4_243;
wire n_0_4_141;
wire n_0_4_142;
wire n_0_4_143;
wire n_0_4_244;
wire n_0_4_145;
wire n_0_4_146;
wire n_0_4_147;
wire n_0_4_148;
wire n_0_4_149;
wire n_0_4_150;
wire n_0_4_151;
wire n_0_4_152;
wire n_0_4_153;
wire n_0_4_154;
wire n_0_4_155;
wire n_0_4_245;
wire n_0_4_157;
wire n_0_4_158;
wire n_0_4_159;
wire n_0_4_246;
wire n_0_4_161;
wire n_0_4_162;
wire n_0_4_163;
wire n_0_4_164;
wire n_0_4_165;
wire n_0_4_166;
wire n_0_4_160;
wire n_0_4_169;
wire n_0_4_170;
wire n_0_4_171;
wire n_0_4_167;
wire n_0_4_173;
wire n_0_4_174;
wire n_0_4_175;
wire n_0_4_176;
wire n_0_4_177;
wire n_0_4_178;
wire n_0_4_179;
wire n_0_4_180;
wire n_0_4_181;
wire n_0_4_182;
wire n_0_4_183;
wire n_0_4_168;
wire n_0_4_185;
wire n_0_4_186;
wire n_0_4_187;
wire n_0_4_172;
wire n_0_4_189;
wire n_0_4_190;
wire n_0_4_191;
wire n_0_4_192;
wire n_0_4_193;
wire n_0_4_194;
wire n_0_4_233;
wire n_0_4_197;
wire n_0_4_198;
wire n_0_4_199;
wire n_0_4_200;
wire n_0_4_201;
wire n_0_4_234;
wire n_0_4_203;
wire n_0_4_204;
wire n_0_4_205;
wire n_0_4_206;
wire n_0_4_207;
wire n_0_4_208;
wire n_0_4_209;
wire n_0_4_210;
wire n_0_4_211;
wire n_0_4_212;
wire n_0_4_213;
wire n_0_4_235;
wire n_0_4_215;
wire n_0_4_216;
wire n_0_4_217;
wire n_0_4_218;
wire n_0_4_220;
wire n_0_4_236;
wire n_0_4_222;
wire n_0_4_223;
wire n_0_4_224;
wire n_0_4_225;
wire n_0_4_226;
wire n_0_4_227;
wire n_0_4_228;
wire n_0_4_231;
wire n_0_4_184;
wire n_0_4_188;
wire n_0_4_195;
wire n_0_4_196;
wire n_0_4_202;
wire n_0_4_214;
wire n_0_4_219;
wire n_0_4_221;
wire n_0_4_229;
wire n_0_4_230;
wire n_0_4_232;
wire n_0_68;
wire n_0_67;
wire n_0_4_237;
wire n_0_4_238;
wire n_0_4_239;
wire n_0_4_240;
wire n_0_4_241;
wire n_0_4_242;
wire n_0_4_247;
wire n_0_4_248;
wire n_0_4_249;
wire n_0_4_250;
wire n_0_4_251;
wire n_0_4_252;
wire n_0_4_257;
wire n_0_4_258;
wire n_0_4_259;
wire n_0_4_260;
wire n_0_4_261;
wire n_0_4_262;
wire sps__n1;
wire sps__n2;
wire sps__n3;
wire sps__n7;
wire sps__n8;
wire sps__n9;
wire sps__n13;
wire sps__n14;
wire sps__n15;
wire sps__n19;
wire sps__n20;
wire sps__n21;
wire sps__n25;
wire sps__n26;
wire sps__n27;
wire sps__n28;
wire sps__n33;
wire sps__n34;
wire sps__n35;
wire sps__n36;
wire sps__n41;
wire sps__n42;
wire sps__n43;
wire sps__n44;
wire sps__n49;
wire sps__n50;
wire sps__n51;
wire sps__n55;
wire sps__n56;
wire sps__n57;
wire sps__n61;
wire sps__n62;
wire sps__n63;
wire sps__n67;
wire sps__n68;
wire sps__n69;
wire sps__n73;
wire sps__n74;
wire sps__n75;
wire sps__n79;
wire sps__n80;
wire sps__n81;
wire sps__n85;
wire sps__n86;
wire sps__n87;
wire sps__n91;
wire sps__n92;
wire sps__n93;
wire sps__n97;
wire sps__n98;
wire sps__n99;
wire sps__n103;
wire sps__n104;
wire sps__n105;
wire sps__n106;
wire sps__n111;
wire sps__n112;
wire sps__n113;
wire sps__n114;
wire sps__n119;
wire sps__n120;
wire sps__n121;
wire sps__n122;
wire sps__n123;

// WARNING . Detected multiport output net(s). Introducing ASSIGN statements.
// This may cause simulation/synthesis mismatches . 
assign doneRead = 1'b1 ;
assign doneWrite = 1'b1 ;

NAND3_X1 i_0_4_270 (.ZN (n_0_4_262), .A1 (n_0_4_260), .A2 (n_0_4_261), .A3 (n_0_5));
NAND2_X1 i_0_4_253 (.ZN (n_0_4_261), .A1 (n_0_4_105), .A2 (n_0_4_109));
NAND2_X1 i_0_4_252 (.ZN (n_0_4_260), .A1 (n_0_4_89), .A2 (n_0_4_93));
NAND3_X1 i_0_4_269 (.ZN (n_0_4_259), .A1 (n_0_4_257), .A2 (n_0_4_258), .A3 (n_0_5));
NAND2_X1 i_0_4_268 (.ZN (n_0_4_258), .A1 (n_0_4_255), .A2 (n_0_4_256));
NAND2_X1 i_0_4_267 (.ZN (n_0_4_257), .A1 (n_0_4_253), .A2 (n_0_4_254));
NAND3_X1 i_0_4_266 (.ZN (n_0_4_252), .A1 (n_0_4_250), .A2 (n_0_4_251), .A3 (n_0_5));
NAND2_X1 i_0_4_265 (.ZN (n_0_4_251), .A1 (n_0_4_144), .A2 (n_0_4_156));
NAND2_X1 i_0_4_264 (.ZN (n_0_4_250), .A1 (n_0_4_139), .A2 (n_0_4_140));
NAND3_X1 i_0_4_263 (.ZN (n_0_4_249), .A1 (n_0_4_247), .A2 (n_0_4_248), .A3 (n_0_5));
NAND2_X1 i_0_4_262 (.ZN (n_0_4_248), .A1 (n_0_4_245), .A2 (n_0_4_246));
NAND2_X1 i_0_4_261 (.ZN (n_0_4_247), .A1 (n_0_4_243), .A2 (n_0_4_244));
NAND3_X1 i_0_4_260 (.ZN (n_0_4_242), .A1 (n_0_4_240), .A2 (n_0_4_241), .A3 (n_0_5));
NAND2_X1 i_0_4_259 (.ZN (n_0_4_241), .A1 (n_0_4_168), .A2 (n_0_4_172));
NAND2_X1 i_0_4_258 (.ZN (n_0_4_240), .A1 (n_0_4_160), .A2 (n_0_4_167));
NAND3_X1 i_0_4_257 (.ZN (n_0_4_239), .A1 (n_0_4_237), .A2 (n_0_4_238), .A3 (n_0_5));
NAND2_X1 i_0_4_256 (.ZN (n_0_4_238), .A1 (n_0_4_235), .A2 (n_0_4_236));
NAND2_X1 i_0_4_255 (.ZN (n_0_4_237), .A1 (n_0_4_233), .A2 (n_0_4_234));
AOI22_X1 i_0_4_254 (.ZN (n_0_67), .A1 (n_0_4_12), .A2 (n_0_4_16), .B1 (n_0_4_32), .B2 (n_0_4_28));
AOI22_X1 i_0_4_251 (.ZN (n_0_68), .A1 (n_0_4_39), .A2 (n_0_4_43), .B1 (n_0_4_59), .B2 (n_0_4_55));
INV_X1 i_0_4_249 (.ZN (n_0_4_232), .A (sps__n103));
NAND3_X1 i_0_4_250 (.ZN (n_0_4_230), .A1 (n_0_4_184), .A2 (\mem[5][0] ), .A3 (sps__n121));
NAND3_X1 i_0_4_243 (.ZN (n_0_4_229), .A1 (n_0_4_184), .A2 (\mem[5][1] ), .A3 (sps__n121));
NAND3_X1 i_0_4_248 (.ZN (n_0_4_221), .A1 (n_0_4_184), .A2 (\mem[5][2] ), .A3 (sps__n121));
NAND3_X1 i_0_4_247 (.ZN (n_0_4_219), .A1 (n_0_4_184), .A2 (\mem[5][3] ), .A3 (sps__n121));
NAND3_X1 i_0_4_246 (.ZN (n_0_4_214), .A1 (n_0_4_184), .A2 (\mem[5][4] ), .A3 (sps__n121));
NAND3_X1 i_0_4_245 (.ZN (n_0_4_202), .A1 (n_0_4_184), .A2 (\mem[5][11] ), .A3 (sps__n121));
NAND3_X1 i_0_4_244 (.ZN (n_0_4_196), .A1 (n_0_4_184), .A2 (\mem[5][13] ), .A3 (sps__n121));
NAND2_X1 i_0_4_240 (.ZN (n_0_4_195), .A1 (n_0_4_184), .A2 (sps__n112));
NAND3_X1 i_0_4_242 (.ZN (n_0_4_188), .A1 (n_0_4_184), .A2 (\mem[5][14] ), .A3 (sps__n121));
INV_X1 i_0_4_241 (.ZN (n_0_4_184), .A (sps__n103));
INV_X2 i_0_4_231 (.ZN (n_0_4_231), .A (sps__n112));
INV_X2 i_0_4_239 (.ZN (n_0_4_228), .A (sps__n121));
INV_X1 i_0_4_238 (.ZN (n_0_4_227), .A (\mem[9][14] ));
NAND2_X1 i_0_4_237 (.ZN (n_0_4_226), .A1 (sps__n106), .A2 (n_0_4_227));
INV_X1 i_0_4_236 (.ZN (n_0_4_225), .A (\mem[1][14] ));
NAND2_X1 i_0_4_235 (.ZN (n_0_4_224), .A1 (n_0_4_232), .A2 (n_0_4_225));
NAND3_X1 i_0_4_234 (.ZN (n_0_4_223), .A1 (n_0_4_224), .A2 (n_0_4_228), .A3 (n_0_4_226));
NAND2_X1 i_0_4_233 (.ZN (n_0_4_222), .A1 (n_0_4_223), .A2 (n_0_4_188));
NAND2_X1 i_0_4_232 (.ZN (n_0_4_236), .A1 (n_0_4_222), .A2 (n_0_4_231));
INV_X1 i_0_4_230 (.ZN (n_0_4_220), .A (sps__n97));
INV_X1 i_0_4_213 (.ZN (n_0_4_218), .A (n_0_4_195));
INV_X1 i_0_4_229 (.ZN (n_0_4_217), .A (\mem[3][14] ));
NAND2_X1 i_0_4_228 (.ZN (n_0_4_216), .A1 (sps__n121), .A2 (\mem[7][14] ));
OAI21_X1 i_0_4_227 (.ZN (n_0_4_215), .A (n_0_4_216), .B1 (n_0_4_217), .B2 (sps__n121));
AOI21_X1 i_0_4_226 (.ZN (n_0_4_235), .A (n_0_4_220), .B1 (n_0_4_215), .B2 (n_0_4_218));
INV_X1 i_0_4_225 (.ZN (n_0_4_213), .A (\mem[6][14] ));
NAND2_X1 i_0_4_224 (.ZN (n_0_4_212), .A1 (address[2]), .A2 (n_0_4_213));
INV_X1 i_0_4_223 (.ZN (n_0_4_211), .A (\mem[2][14] ));
NAND2_X1 i_0_4_222 (.ZN (n_0_4_210), .A1 (n_0_4_228), .A2 (n_0_4_211));
NAND3_X1 i_0_4_221 (.ZN (n_0_4_209), .A1 (n_0_4_210), .A2 (sps__n113), .A3 (n_0_4_212));
INV_X1 i_0_4_220 (.ZN (n_0_4_208), .A (\mem[4][14] ));
NAND2_X1 i_0_4_219 (.ZN (n_0_4_207), .A1 (address[2]), .A2 (n_0_4_208));
INV_X1 i_0_4_218 (.ZN (n_0_4_206), .A (\mem[0][14] ));
NAND2_X1 i_0_4_217 (.ZN (n_0_4_205), .A1 (n_0_4_228), .A2 (n_0_4_206));
NAND3_X1 i_0_4_216 (.ZN (n_0_4_204), .A1 (n_0_4_205), .A2 (n_0_4_231), .A3 (n_0_4_207));
NAND2_X1 i_0_4_215 (.ZN (n_0_4_203), .A1 (n_0_4_209), .A2 (n_0_4_204));
NAND2_X1 i_0_4_214 (.ZN (n_0_4_234), .A1 (n_0_4_203), .A2 (n_0_4_232));
NAND2_X1 i_0_4_212 (.ZN (n_0_4_201), .A1 (n_0_4_228), .A2 (sps__n103));
INV_X1 i_0_4_68 (.ZN (n_0_4_200), .A (n_0_4_201));
INV_X1 i_0_4_211 (.ZN (n_0_4_199), .A (\mem[8][14] ));
NAND2_X1 i_0_4_210 (.ZN (n_0_4_198), .A1 (sps__n113), .A2 (\mem[10][14] ));
OAI21_X1 i_0_4_209 (.ZN (n_0_4_197), .A (n_0_4_198), .B1 (n_0_4_199), .B2 (sps__n113));
AOI21_X1 i_0_4_208 (.ZN (n_0_4_233), .A (sps__n97), .B1 (n_0_4_197), .B2 (n_0_4_200));
INV_X1 i_0_4_207 (.ZN (n_0_4_194), .A (\mem[9][13] ));
NAND2_X1 i_0_4_206 (.ZN (n_0_4_193), .A1 (sps__n103), .A2 (n_0_4_194));
INV_X1 i_0_4_205 (.ZN (n_0_4_192), .A (\mem[1][13] ));
NAND2_X1 i_0_4_204 (.ZN (n_0_4_191), .A1 (n_0_4_232), .A2 (n_0_4_192));
NAND3_X1 i_0_4_203 (.ZN (n_0_4_190), .A1 (n_0_4_191), .A2 (n_0_4_228), .A3 (n_0_4_193));
NAND2_X1 i_0_4_202 (.ZN (n_0_4_189), .A1 (n_0_4_190), .A2 (n_0_4_196));
NAND2_X1 i_0_4_201 (.ZN (n_0_4_172), .A1 (n_0_4_189), .A2 (n_0_4_231));
INV_X1 i_0_4_200 (.ZN (n_0_4_187), .A (\mem[3][13] ));
NAND2_X1 i_0_4_199 (.ZN (n_0_4_186), .A1 (sps__n121), .A2 (\mem[7][13] ));
OAI21_X1 i_0_4_198 (.ZN (n_0_4_185), .A (n_0_4_186), .B1 (n_0_4_187), .B2 (sps__n121));
AOI21_X1 i_0_4_197 (.ZN (n_0_4_168), .A (n_0_4_220), .B1 (n_0_4_185), .B2 (n_0_4_218));
INV_X1 i_0_4_196 (.ZN (n_0_4_183), .A (\mem[6][13] ));
NAND2_X1 i_0_4_195 (.ZN (n_0_4_182), .A1 (sps__n121), .A2 (n_0_4_183));
INV_X1 i_0_4_194 (.ZN (n_0_4_181), .A (\mem[2][13] ));
NAND2_X1 i_0_4_193 (.ZN (n_0_4_180), .A1 (n_0_4_228), .A2 (n_0_4_181));
NAND3_X1 i_0_4_192 (.ZN (n_0_4_179), .A1 (n_0_4_180), .A2 (sps__n112), .A3 (n_0_4_182));
INV_X1 i_0_4_191 (.ZN (n_0_4_178), .A (\mem[4][13] ));
NAND2_X1 i_0_4_190 (.ZN (n_0_4_177), .A1 (sps__n121), .A2 (n_0_4_178));
INV_X1 i_0_4_189 (.ZN (n_0_4_176), .A (\mem[0][13] ));
NAND2_X1 i_0_4_188 (.ZN (n_0_4_175), .A1 (n_0_4_228), .A2 (n_0_4_176));
NAND3_X1 i_0_4_187 (.ZN (n_0_4_174), .A1 (n_0_4_175), .A2 (n_0_4_231), .A3 (n_0_4_177));
NAND2_X1 i_0_4_186 (.ZN (n_0_4_173), .A1 (n_0_4_179), .A2 (n_0_4_174));
NAND2_X1 i_0_4_185 (.ZN (n_0_4_167), .A1 (n_0_4_173), .A2 (n_0_4_232));
INV_X1 i_0_4_184 (.ZN (n_0_4_171), .A (\mem[8][13] ));
NAND2_X1 i_0_4_183 (.ZN (n_0_4_170), .A1 (sps__n112), .A2 (\mem[10][13] ));
OAI21_X1 i_0_4_182 (.ZN (n_0_4_169), .A (n_0_4_170), .B1 (n_0_4_171), .B2 (sps__n112));
AOI21_X1 i_0_4_181 (.ZN (n_0_4_160), .A (sps__n99), .B1 (n_0_4_169), .B2 (n_0_4_200));
INV_X1 i_0_4_180 (.ZN (n_0_4_166), .A (\mem[9][11] ));
NAND2_X1 i_0_4_179 (.ZN (n_0_4_165), .A1 (sps__n103), .A2 (n_0_4_166));
INV_X1 i_0_4_178 (.ZN (n_0_4_164), .A (\mem[1][11] ));
NAND2_X1 i_0_4_177 (.ZN (n_0_4_163), .A1 (n_0_4_232), .A2 (n_0_4_164));
NAND3_X1 i_0_4_176 (.ZN (n_0_4_162), .A1 (n_0_4_163), .A2 (n_0_4_228), .A3 (n_0_4_165));
NAND2_X1 i_0_4_175 (.ZN (n_0_4_161), .A1 (n_0_4_162), .A2 (n_0_4_202));
NAND2_X1 i_0_4_174 (.ZN (n_0_4_246), .A1 (n_0_4_161), .A2 (n_0_4_231));
INV_X1 i_0_4_173 (.ZN (n_0_4_159), .A (\mem[3][11] ));
NAND2_X1 i_0_4_172 (.ZN (n_0_4_158), .A1 (sps__n121), .A2 (\mem[7][11] ));
OAI21_X1 i_0_4_171 (.ZN (n_0_4_157), .A (n_0_4_158), .B1 (n_0_4_159), .B2 (sps__n121));
AOI21_X1 i_0_4_170 (.ZN (n_0_4_245), .A (n_0_4_220), .B1 (n_0_4_157), .B2 (n_0_4_218));
INV_X1 i_0_4_169 (.ZN (n_0_4_155), .A (\mem[6][11] ));
NAND2_X1 i_0_4_168 (.ZN (n_0_4_154), .A1 (sps__n121), .A2 (n_0_4_155));
INV_X1 i_0_4_167 (.ZN (n_0_4_153), .A (\mem[2][11] ));
NAND2_X1 i_0_4_166 (.ZN (n_0_4_152), .A1 (n_0_4_228), .A2 (n_0_4_153));
NAND3_X1 i_0_4_165 (.ZN (n_0_4_151), .A1 (n_0_4_152), .A2 (sps__n112), .A3 (n_0_4_154));
INV_X1 i_0_4_164 (.ZN (n_0_4_150), .A (\mem[4][11] ));
NAND2_X1 i_0_4_163 (.ZN (n_0_4_149), .A1 (sps__n121), .A2 (n_0_4_150));
INV_X1 i_0_4_162 (.ZN (n_0_4_148), .A (\mem[0][11] ));
NAND2_X1 i_0_4_161 (.ZN (n_0_4_147), .A1 (n_0_4_228), .A2 (n_0_4_148));
NAND3_X1 i_0_4_160 (.ZN (n_0_4_146), .A1 (n_0_4_147), .A2 (n_0_4_231), .A3 (n_0_4_149));
NAND2_X1 i_0_4_159 (.ZN (n_0_4_145), .A1 (n_0_4_151), .A2 (n_0_4_146));
NAND2_X1 i_0_4_158 (.ZN (n_0_4_244), .A1 (n_0_4_145), .A2 (n_0_4_232));
INV_X1 i_0_4_157 (.ZN (n_0_4_143), .A (\mem[8][11] ));
NAND2_X1 i_0_4_156 (.ZN (n_0_4_142), .A1 (sps__n112), .A2 (\mem[10][11] ));
OAI21_X1 i_0_4_155 (.ZN (n_0_4_141), .A (n_0_4_142), .B1 (n_0_4_143), .B2 (sps__n112));
AOI21_X1 i_0_4_154 (.ZN (n_0_4_243), .A (sps__n99), .B1 (n_0_4_141), .B2 (n_0_4_200));
INV_X1 i_0_4_153 (.ZN (n_0_4_138), .A (\mem[9][4] ));
NAND2_X1 i_0_4_152 (.ZN (n_0_4_137), .A1 (sps__n103), .A2 (n_0_4_138));
INV_X1 i_0_4_151 (.ZN (n_0_4_136), .A (\mem[1][4] ));
NAND2_X1 i_0_4_150 (.ZN (n_0_4_135), .A1 (n_0_4_232), .A2 (n_0_4_136));
NAND3_X1 i_0_4_149 (.ZN (n_0_4_134), .A1 (n_0_4_135), .A2 (n_0_4_228), .A3 (n_0_4_137));
NAND2_X1 i_0_4_148 (.ZN (n_0_4_133), .A1 (n_0_4_134), .A2 (n_0_4_214));
NAND2_X1 i_0_4_147 (.ZN (n_0_4_156), .A1 (n_0_4_133), .A2 (n_0_4_231));
INV_X1 i_0_4_146 (.ZN (n_0_4_132), .A (\mem[3][4] ));
NAND2_X1 i_0_4_145 (.ZN (n_0_4_131), .A1 (sps__n121), .A2 (\mem[7][4] ));
OAI21_X1 i_0_4_144 (.ZN (n_0_4_130), .A (n_0_4_131), .B1 (n_0_4_132), .B2 (sps__n121));
AOI21_X1 i_0_4_143 (.ZN (n_0_4_144), .A (n_0_4_220), .B1 (n_0_4_130), .B2 (n_0_4_218));
INV_X1 i_0_4_142 (.ZN (n_0_4_129), .A (\mem[6][4] ));
NAND2_X1 i_0_4_141 (.ZN (n_0_4_128), .A1 (sps__n122), .A2 (n_0_4_129));
INV_X1 i_0_4_140 (.ZN (n_0_4_127), .A (\mem[2][4] ));
NAND2_X1 i_0_4_139 (.ZN (n_0_4_126), .A1 (n_0_4_228), .A2 (n_0_4_127));
NAND3_X1 i_0_4_138 (.ZN (n_0_4_125), .A1 (n_0_4_126), .A2 (sps__n112), .A3 (n_0_4_128));
INV_X1 i_0_4_137 (.ZN (n_0_4_124), .A (\mem[4][4] ));
NAND2_X1 i_0_4_136 (.ZN (n_0_4_123), .A1 (sps__n122), .A2 (n_0_4_124));
INV_X1 i_0_4_135 (.ZN (n_0_4_122), .A (\mem[0][4] ));
NAND2_X1 i_0_4_134 (.ZN (n_0_4_121), .A1 (n_0_4_228), .A2 (n_0_4_122));
NAND3_X1 i_0_4_133 (.ZN (n_0_4_120), .A1 (n_0_4_121), .A2 (n_0_4_231), .A3 (n_0_4_123));
NAND2_X1 i_0_4_132 (.ZN (n_0_4_119), .A1 (n_0_4_125), .A2 (n_0_4_120));
NAND2_X1 i_0_4_131 (.ZN (n_0_4_140), .A1 (n_0_4_119), .A2 (n_0_4_232));
INV_X1 i_0_4_130 (.ZN (n_0_4_118), .A (\mem[8][4] ));
NAND2_X1 i_0_4_129 (.ZN (n_0_4_117), .A1 (sps__n112), .A2 (\mem[10][4] ));
OAI21_X1 i_0_4_128 (.ZN (n_0_4_116), .A (n_0_4_117), .B1 (n_0_4_118), .B2 (sps__n112));
AOI21_X1 i_0_4_127 (.ZN (n_0_4_139), .A (sps__n99), .B1 (n_0_4_116), .B2 (n_0_4_200));
INV_X1 i_0_4_126 (.ZN (n_0_4_115), .A (\mem[9][3] ));
NAND2_X1 i_0_4_125 (.ZN (n_0_4_114), .A1 (sps__n104), .A2 (n_0_4_115));
INV_X1 i_0_4_124 (.ZN (n_0_4_113), .A (\mem[1][3] ));
NAND2_X1 i_0_4_123 (.ZN (n_0_4_112), .A1 (n_0_4_232), .A2 (n_0_4_113));
NAND3_X1 i_0_4_122 (.ZN (n_0_4_111), .A1 (n_0_4_112), .A2 (n_0_4_228), .A3 (n_0_4_114));
NAND2_X1 i_0_4_121 (.ZN (n_0_4_110), .A1 (n_0_4_111), .A2 (n_0_4_219));
NAND2_X1 i_0_4_120 (.ZN (n_0_4_256), .A1 (n_0_4_110), .A2 (n_0_4_231));
INV_X1 i_0_4_119 (.ZN (n_0_4_108), .A (\mem[3][3] ));
NAND2_X1 i_0_4_118 (.ZN (n_0_4_107), .A1 (sps__n121), .A2 (\mem[7][3] ));
OAI21_X1 i_0_4_117 (.ZN (n_0_4_106), .A (n_0_4_107), .B1 (n_0_4_108), .B2 (sps__n121));
AOI21_X1 i_0_4_116 (.ZN (n_0_4_255), .A (n_0_4_220), .B1 (n_0_4_106), .B2 (n_0_4_218));
INV_X1 i_0_4_115 (.ZN (n_0_4_104), .A (\mem[6][3] ));
NAND2_X1 i_0_4_114 (.ZN (n_0_4_103), .A1 (sps__n122), .A2 (n_0_4_104));
INV_X1 i_0_4_113 (.ZN (n_0_4_102), .A (\mem[2][3] ));
NAND2_X1 i_0_4_112 (.ZN (n_0_4_101), .A1 (n_0_4_228), .A2 (n_0_4_102));
NAND3_X1 i_0_4_111 (.ZN (n_0_4_100), .A1 (n_0_4_101), .A2 (sps__n112), .A3 (n_0_4_103));
INV_X1 i_0_4_110 (.ZN (n_0_4_99), .A (\mem[4][3] ));
NAND2_X1 i_0_4_109 (.ZN (n_0_4_98), .A1 (sps__n122), .A2 (n_0_4_99));
INV_X1 i_0_4_108 (.ZN (n_0_4_97), .A (\mem[0][3] ));
NAND2_X1 i_0_4_107 (.ZN (n_0_4_96), .A1 (n_0_4_228), .A2 (n_0_4_97));
NAND3_X1 i_0_4_106 (.ZN (n_0_4_95), .A1 (n_0_4_96), .A2 (n_0_4_231), .A3 (n_0_4_98));
NAND2_X1 i_0_4_105 (.ZN (n_0_4_94), .A1 (n_0_4_100), .A2 (n_0_4_95));
NAND2_X1 i_0_4_104 (.ZN (n_0_4_254), .A1 (n_0_4_94), .A2 (n_0_4_232));
INV_X1 i_0_4_103 (.ZN (n_0_4_92), .A (\mem[8][3] ));
NAND2_X1 i_0_4_102 (.ZN (n_0_4_91), .A1 (sps__n112), .A2 (\mem[10][3] ));
OAI21_X1 i_0_4_101 (.ZN (n_0_4_90), .A (n_0_4_91), .B1 (n_0_4_92), .B2 (sps__n112));
AOI21_X1 i_0_4_100 (.ZN (n_0_4_253), .A (sps__n99), .B1 (n_0_4_90), .B2 (n_0_4_200));
INV_X1 i_0_4_99 (.ZN (n_0_4_88), .A (\mem[9][2] ));
NAND2_X1 i_0_4_98 (.ZN (n_0_4_87), .A1 (sps__n103), .A2 (n_0_4_88));
INV_X1 i_0_4_97 (.ZN (n_0_4_86), .A (\mem[1][2] ));
NAND2_X1 i_0_4_96 (.ZN (n_0_4_85), .A1 (n_0_4_232), .A2 (n_0_4_86));
NAND3_X1 i_0_4_95 (.ZN (n_0_4_84), .A1 (n_0_4_85), .A2 (n_0_4_228), .A3 (n_0_4_87));
NAND2_X1 i_0_4_94 (.ZN (n_0_4_83), .A1 (n_0_4_84), .A2 (n_0_4_221));
NAND2_X1 i_0_4_93 (.ZN (n_0_4_109), .A1 (n_0_4_83), .A2 (n_0_4_231));
INV_X1 i_0_4_92 (.ZN (n_0_4_82), .A (\mem[3][2] ));
NAND2_X1 i_0_4_91 (.ZN (n_0_4_81), .A1 (sps__n121), .A2 (\mem[7][2] ));
OAI21_X1 i_0_4_90 (.ZN (n_0_4_80), .A (n_0_4_81), .B1 (n_0_4_82), .B2 (sps__n121));
AOI21_X1 i_0_4_89 (.ZN (n_0_4_105), .A (n_0_4_220), .B1 (n_0_4_80), .B2 (n_0_4_218));
INV_X1 i_0_4_88 (.ZN (n_0_4_79), .A (\mem[6][2] ));
NAND2_X1 i_0_4_87 (.ZN (n_0_4_78), .A1 (sps__n121), .A2 (n_0_4_79));
INV_X1 i_0_4_86 (.ZN (n_0_4_77), .A (\mem[2][2] ));
NAND2_X1 i_0_4_85 (.ZN (n_0_4_76), .A1 (n_0_4_228), .A2 (n_0_4_77));
NAND3_X1 i_0_4_84 (.ZN (n_0_4_75), .A1 (n_0_4_76), .A2 (sps__n112), .A3 (n_0_4_78));
INV_X1 i_0_4_83 (.ZN (n_0_4_74), .A (\mem[4][2] ));
NAND2_X1 i_0_4_82 (.ZN (n_0_4_73), .A1 (sps__n121), .A2 (n_0_4_74));
INV_X1 i_0_4_81 (.ZN (n_0_4_72), .A (\mem[0][2] ));
NAND2_X1 i_0_4_80 (.ZN (n_0_4_71), .A1 (n_0_4_228), .A2 (n_0_4_72));
NAND3_X1 i_0_4_79 (.ZN (n_0_4_70), .A1 (n_0_4_71), .A2 (n_0_4_231), .A3 (n_0_4_73));
NAND2_X1 i_0_4_78 (.ZN (n_0_4_69), .A1 (n_0_4_75), .A2 (n_0_4_70));
NAND2_X1 i_0_4_77 (.ZN (n_0_4_93), .A1 (n_0_4_69), .A2 (n_0_4_232));
INV_X1 i_0_4_76 (.ZN (n_0_4_68), .A (\mem[8][2] ));
NAND2_X1 i_0_4_75 (.ZN (n_0_4_67), .A1 (sps__n112), .A2 (\mem[10][2] ));
OAI21_X1 i_0_4_74 (.ZN (n_0_4_66), .A (n_0_4_67), .B1 (n_0_4_68), .B2 (sps__n112));
AOI21_X1 i_0_4_73 (.ZN (n_0_4_89), .A (sps__n97), .B1 (n_0_4_66), .B2 (n_0_4_200));
INV_X1 i_0_4_72 (.ZN (n_0_4_65), .A (\mem[9][1] ));
NAND2_X1 i_0_4_71 (.ZN (n_0_4_64), .A1 (sps__n103), .A2 (n_0_4_65));
INV_X1 i_0_4_70 (.ZN (n_0_4_63), .A (\mem[1][1] ));
NAND2_X1 i_0_4_69 (.ZN (n_0_4_62), .A1 (n_0_4_232), .A2 (n_0_4_63));
NAND3_X1 i_0_4_67 (.ZN (n_0_4_61), .A1 (n_0_4_62), .A2 (n_0_4_228), .A3 (n_0_4_64));
NAND2_X1 i_0_4_66 (.ZN (n_0_4_60), .A1 (n_0_4_61), .A2 (n_0_4_229));
NAND2_X1 i_0_4_64 (.ZN (n_0_4_59), .A1 (n_0_4_60), .A2 (n_0_4_231));
INV_X1 i_0_4_65 (.ZN (n_0_4_58), .A (\mem[3][1] ));
NAND2_X1 i_0_4_63 (.ZN (n_0_4_57), .A1 (sps__n119), .A2 (\mem[7][1] ));
OAI21_X1 i_0_4_62 (.ZN (n_0_4_56), .A (n_0_4_57), .B1 (n_0_4_58), .B2 (sps__n119));
AOI21_X1 i_0_4_57 (.ZN (n_0_4_55), .A (n_0_4_220), .B1 (n_0_4_56), .B2 (n_0_4_218));
INV_X1 i_0_4_61 (.ZN (n_0_4_54), .A (\mem[6][1] ));
NAND2_X1 i_0_4_60 (.ZN (n_0_4_53), .A1 (sps__n119), .A2 (n_0_4_54));
INV_X1 i_0_4_59 (.ZN (n_0_4_52), .A (\mem[2][1] ));
NAND2_X1 i_0_4_58 (.ZN (n_0_4_51), .A1 (n_0_4_228), .A2 (n_0_4_52));
NAND3_X1 i_0_4_52 (.ZN (n_0_4_50), .A1 (n_0_4_51), .A2 (sps__n113), .A3 (n_0_4_53));
INV_X1 i_0_4_56 (.ZN (n_0_4_49), .A (\mem[4][1] ));
NAND2_X1 i_0_4_55 (.ZN (n_0_4_48), .A1 (sps__n119), .A2 (n_0_4_49));
INV_X1 i_0_4_54 (.ZN (n_0_4_47), .A (\mem[0][1] ));
NAND2_X1 i_0_4_53 (.ZN (n_0_4_46), .A1 (n_0_4_228), .A2 (n_0_4_47));
NAND3_X1 i_0_4_51 (.ZN (n_0_4_45), .A1 (n_0_4_46), .A2 (n_0_4_231), .A3 (n_0_4_48));
NAND2_X1 i_0_4_50 (.ZN (n_0_4_44), .A1 (n_0_4_50), .A2 (n_0_4_45));
NAND2_X1 i_0_4_48 (.ZN (n_0_4_43), .A1 (n_0_4_44), .A2 (n_0_4_232));
INV_X1 i_0_4_49 (.ZN (n_0_4_42), .A (\mem[8][1] ));
NAND2_X1 i_0_4_47 (.ZN (n_0_4_41), .A1 (sps__n113), .A2 (\mem[10][1] ));
OAI21_X1 i_0_4_46 (.ZN (n_0_4_40), .A (n_0_4_41), .B1 (n_0_4_42), .B2 (sps__n113));
AOI21_X1 i_0_4_3 (.ZN (n_0_4_39), .A (sps__n97), .B1 (n_0_4_40), .B2 (n_0_4_200));
INV_X1 i_0_4_45 (.ZN (n_0_4_38), .A (\mem[9][0] ));
NAND2_X1 i_0_4_44 (.ZN (n_0_4_37), .A1 (sps__n106), .A2 (n_0_4_38));
INV_X1 i_0_4_43 (.ZN (n_0_4_36), .A (\mem[1][0] ));
NAND2_X1 i_0_4_42 (.ZN (n_0_4_35), .A1 (n_0_4_232), .A2 (n_0_4_36));
NAND3_X1 i_0_4_41 (.ZN (n_0_4_34), .A1 (n_0_4_35), .A2 (n_0_4_228), .A3 (n_0_4_37));
NAND2_X1 i_0_4_40 (.ZN (n_0_4_33), .A1 (n_0_4_34), .A2 (n_0_4_230));
NAND2_X1 i_0_4_39 (.ZN (n_0_4_32), .A1 (n_0_4_33), .A2 (n_0_4_231));
INV_X1 i_0_4_38 (.ZN (n_0_4_31), .A (\mem[3][0] ));
NAND2_X1 i_0_4_37 (.ZN (n_0_4_30), .A1 (sps__n119), .A2 (\mem[7][0] ));
OAI21_X1 i_0_4_36 (.ZN (n_0_4_29), .A (n_0_4_30), .B1 (n_0_4_31), .B2 (sps__n119));
AOI21_X1 i_0_4_35 (.ZN (n_0_4_28), .A (n_0_4_220), .B1 (n_0_4_29), .B2 (n_0_4_218));
INV_X1 i_0_4_34 (.ZN (n_0_4_27), .A (\mem[6][0] ));
NAND2_X1 i_0_4_33 (.ZN (n_0_4_26), .A1 (sps__n119), .A2 (n_0_4_27));
INV_X1 i_0_4_32 (.ZN (n_0_4_25), .A (\mem[2][0] ));
NAND2_X1 i_0_4_31 (.ZN (n_0_4_24), .A1 (n_0_4_228), .A2 (n_0_4_25));
NAND3_X1 i_0_4_30 (.ZN (n_0_4_23), .A1 (n_0_4_24), .A2 (sps__n113), .A3 (n_0_4_26));
INV_X1 i_0_4_29 (.ZN (n_0_4_22), .A (\mem[4][0] ));
NAND2_X1 i_0_4_28 (.ZN (n_0_4_21), .A1 (sps__n119), .A2 (n_0_4_22));
INV_X1 i_0_4_27 (.ZN (n_0_4_20), .A (\mem[0][0] ));
NAND2_X1 i_0_4_26 (.ZN (n_0_4_19), .A1 (n_0_4_228), .A2 (n_0_4_20));
NAND3_X1 i_0_4_25 (.ZN (n_0_4_18), .A1 (n_0_4_19), .A2 (n_0_4_231), .A3 (n_0_4_21));
NAND2_X1 i_0_4_24 (.ZN (n_0_4_17), .A1 (n_0_4_23), .A2 (n_0_4_18));
NAND2_X1 i_0_4_23 (.ZN (n_0_4_16), .A1 (n_0_4_17), .A2 (n_0_4_232));
INV_X1 i_0_4_22 (.ZN (n_0_4_15), .A (\mem[8][0] ));
NAND2_X1 i_0_4_21 (.ZN (n_0_4_14), .A1 (sps__n113), .A2 (\mem[10][0] ));
OAI21_X1 i_0_4_20 (.ZN (n_0_4_13), .A (n_0_4_14), .B1 (n_0_4_15), .B2 (sps__n113));
AOI21_X1 i_0_4_19 (.ZN (n_0_4_12), .A (sps__n97), .B1 (n_0_4_13), .B2 (n_0_4_200));
INV_X1 i_0_4_18 (.ZN (n_0_4_11), .A (n_0_5));
NAND2_X1 i_0_4_17 (.ZN (n_0_4_10), .A1 (n_0_4_11), .A2 (dataout[14]));
NAND2_X1 i_0_4_16 (.ZN (n_0_8), .A1 (n_0_4_239), .A2 (n_0_4_10));
INV_X1 i_0_4_15 (.ZN (n_0_4_9), .A (n_0_5));
NAND2_X1 i_0_4_14 (.ZN (n_0_4_8), .A1 (n_0_4_9), .A2 (dataout[13]));
NAND2_X1 i_0_4_13 (.ZN (n_0_74), .A1 (n_0_4_242), .A2 (n_0_4_8));
INV_X1 i_0_4_12 (.ZN (n_0_4_7), .A (n_0_5));
NAND2_X1 i_0_4_11 (.ZN (n_0_4_6), .A1 (n_0_4_7), .A2 (dataout[11]));
NAND2_X1 i_0_4_10 (.ZN (n_0_9), .A1 (n_0_4_249), .A2 (n_0_4_6));
INV_X1 i_0_4_9 (.ZN (n_0_4_5), .A (n_0_5));
NAND2_X1 i_0_4_8 (.ZN (n_0_4_4), .A1 (n_0_4_5), .A2 (dataout[4]));
NAND2_X1 i_0_4_7 (.ZN (n_0_73), .A1 (n_0_4_252), .A2 (n_0_4_4));
INV_X1 i_0_4_6 (.ZN (n_0_4_3), .A (n_0_5));
NAND2_X1 i_0_4_5 (.ZN (n_0_4_2), .A1 (n_0_4_3), .A2 (dataout[3]));
NAND2_X1 i_0_4_4 (.ZN (n_0_11), .A1 (n_0_4_259), .A2 (n_0_4_2));
INV_X1 i_0_4_2 (.ZN (n_0_4_1), .A (n_0_5));
NAND2_X1 i_0_4_1 (.ZN (n_0_4_0), .A1 (n_0_4_1), .A2 (dataout[2]));
NAND2_X1 i_0_4_0 (.ZN (n_0_72), .A1 (n_0_4_262), .A2 (n_0_4_0));
DFF_X2 \temp_reg[7]  (.Q (dataout[7]), .CK (n_0_32), .D (n_0_48));
DFF_X2 \temp_reg[8]  (.Q (dataout[8]), .CK (n_0_32), .D (n_0_70));
DFF_X2 \temp_reg[12]  (.Q (dataout[12]), .CK (n_0_32), .D (n_0_71));
DFF_X2 \temp_reg[15]  (.Q (dataout[15]), .CK (n_0_32), .D (n_0_69));
DFF_X1 \temp_reg[0]  (.Q (dataout[0]), .CK (n_0_32), .D (n_0_31));
DFF_X1 \temp_reg[1]  (.Q (dataout[1]), .CK (n_0_32), .D (n_0_13));
DFF_X1 \temp_reg[2]  (.Q (dataout[2]), .CK (n_0_32), .D (n_0_72));
DFF_X1 \temp_reg[3]  (.Q (dataout[3]), .CK (n_0_32), .D (n_0_11));
DFF_X1 \temp_reg[4]  (.Q (dataout[4]), .CK (n_0_32), .D (n_0_73));
DFF_X1 \temp_reg[11]  (.Q (dataout[11]), .CK (n_0_32), .D (n_0_9));
DFF_X1 \temp_reg[13]  (.Q (dataout[13]), .CK (n_0_32), .D (n_0_74));
DFF_X1 \temp_reg[14]  (.Q (dataout[14]), .CK (n_0_32), .D (n_0_8));
NAND3_X1 i_0_1_37 (.ZN (n_0_7), .A1 (n_0_1_34), .A2 (n_0_1_35), .A3 (n_0_1_36));
NAND2_X1 i_0_1_36 (.ZN (n_0_1_36), .A1 (n_0_1_25), .A2 (\mem[0][0] ));
NAND3_X1 i_0_1_35 (.ZN (n_0_1_35), .A1 (n_0_1_27), .A2 (n_0_1_33), .A3 (n_0_1_30));
NAND2_X1 i_0_1_34 (.ZN (n_0_1_34), .A1 (n_0_1_24), .A2 (\mem[0][0] ));
NOR2_X1 i_0_1_33 (.ZN (n_0_1_33), .A1 (n_0_1_0), .A2 (n_0_1_19));
INV_X1 i_0_1_32 (.ZN (n_0_1_32), .A (n_0_1_19));
INV_X1 i_0_1_31 (.ZN (n_0_1_31), .A (n_0_1_0));
NOR2_X1 i_0_1_30 (.ZN (n_0_1_30), .A1 (n_0_1_5), .A2 (n_0_1_15));
INV_X1 i_0_1_29 (.ZN (n_0_1_29), .A (n_0_1_15));
INV_X1 i_0_1_28 (.ZN (n_0_1_28), .A (n_0_1_5));
INV_X1 i_0_1_27 (.ZN (n_0_1_27), .A (n_0_1_26));
NAND2_X1 i_0_1_26 (.ZN (n_0_1_26), .A1 (n_0_1_10), .A2 (data[0]));
NAND2_X1 i_0_1_25 (.ZN (n_0_1_25), .A1 (n_0_1_31), .A2 (n_0_1_28));
NAND3_X1 i_0_1_24 (.ZN (n_0_1_24), .A1 (n_0_1_32), .A2 (n_0_1_29), .A3 (n_0_1_10));
INV_X1 i_0_1_23 (.ZN (n_0_1_23), .A (sps__n35));
INV_X1 i_0_1_22 (.ZN (n_0_1_22), .A (sps__n8));
INV_X1 i_0_1_21 (.ZN (n_0_1_21), .A (sps__n13));
INV_X1 i_0_1_20 (.ZN (n_0_1_20), .A (sps__n49));
NAND4_X1 i_0_1_19 (.ZN (n_0_1_19), .A1 (n_0_1_23), .A2 (n_0_1_22), .A3 (n_0_1_21), .A4 (n_0_1_20));
INV_X1 i_0_1_18 (.ZN (n_0_1_18), .A (sps__n61));
INV_X1 i_0_1_17 (.ZN (n_0_1_17), .A (sps__n73));
INV_X1 i_0_1_12 (.ZN (n_0_1_16), .A (sps__n85));
NAND4_X1 i_0_1_11 (.ZN (n_0_1_15), .A1 (n_0_1_18), .A2 (n_0_1_17), .A3 (n_0_1_16), .A4 (sps__n1));
INV_X1 i_0_1_6 (.ZN (n_0_1_14), .A (sps__n119));
INV_X1 i_0_1_5 (.ZN (n_0_1_13), .A (sps__n112));
INV_X1 i_0_1_4 (.ZN (n_0_1_12), .A (sps__n97));
NAND3_X1 i_0_1_1 (.ZN (n_0_1_11), .A1 (n_0_1_14), .A2 (n_0_1_13), .A3 (n_0_1_12));
INV_X1 i_0_1_0 (.ZN (n_0_1_10), .A (n_0_1_11));
INV_X1 i_0_1_16 (.ZN (n_0_1_9), .A (sps__n67));
INV_X1 i_0_1_15 (.ZN (n_0_1_8), .A (sps__n21));
INV_X1 i_0_1_14 (.ZN (n_0_1_7), .A (sps__n79));
INV_X1 i_0_1_13 (.ZN (n_0_1_6), .A (sps__n106));
NAND4_X1 i_0_1_3 (.ZN (n_0_1_5), .A1 (n_0_1_9), .A2 (n_0_1_8), .A3 (n_0_1_7), .A4 (n_0_1_6));
INV_X1 i_0_1_10 (.ZN (n_0_1_4), .A (sps__n56));
INV_X1 i_0_1_9 (.ZN (n_0_1_3), .A (sps__n27));
INV_X1 i_0_1_8 (.ZN (n_0_1_2), .A (sps__n41));
INV_X1 i_0_1_7 (.ZN (n_0_1_1), .A (sps__n93));
NAND4_X1 i_0_1_2 (.ZN (n_0_1_0), .A1 (n_0_1_4), .A2 (n_0_1_3), .A3 (n_0_1_2), .A4 (n_0_1_1));
OAI21_X1 i_0_189_6 (.ZN (n_0_189_35), .A (\mem[8][0] ), .B1 (n_0_189_10), .B2 (n_0_189_14));
NAND4_X1 i_0_189_28 (.ZN (n_0_189_34), .A1 (n_0_189_9), .A2 (n_0_189_7), .A3 (n_0_189_8), .A4 (data[0]));
NAND2_X1 i_0_189_27 (.ZN (n_0_189_33), .A1 (n_0_189_32), .A2 (\mem[8][0] ));
NAND3_X1 i_0_189_38 (.ZN (n_0_189_32), .A1 (n_0_189_29), .A2 (n_0_189_30), .A3 (n_0_189_31));
INV_X1 i_0_189_37 (.ZN (n_0_189_31), .A (n_0_189_24));
INV_X1 i_0_189_36 (.ZN (n_0_189_30), .A (n_0_189_25));
NOR2_X1 i_0_189_29 (.ZN (n_0_189_29), .A1 (n_0_189_23), .A2 (n_0_189_26));
NAND3_X1 i_0_189_26 (.ZN (n_0_6), .A1 (n_0_189_28), .A2 (n_0_189_33), .A3 (n_0_189_35));
NAND3_X1 i_0_189_23 (.ZN (n_0_189_28), .A1 (n_0_189_19), .A2 (n_0_189_27), .A3 (n_0_189_20));
NOR2_X1 i_0_189_24 (.ZN (n_0_189_27), .A1 (n_0_189_14), .A2 (n_0_189_22));
NAND2_X1 i_0_189_44 (.ZN (n_0_189_26), .A1 (n_0_189_7), .A2 (n_0_189_8));
NAND3_X1 i_0_189_5 (.ZN (n_0_189_25), .A1 (n_0_189_3), .A2 (n_0_189_6), .A3 (sps__n106));
NAND3_X1 i_0_189_40 (.ZN (n_0_189_24), .A1 (n_0_189_0), .A2 (n_0_189_9), .A3 (n_0_189_1));
NAND3_X1 i_0_189_35 (.ZN (n_0_189_23), .A1 (n_0_189_4), .A2 (n_0_189_2), .A3 (n_0_189_5));
NAND4_X1 i_0_189_22 (.ZN (n_0_189_22), .A1 (n_0_189_3), .A2 (n_0_189_2), .A3 (n_0_189_1), .A4 (n_0_189_0));
NAND4_X1 i_0_189_17 (.ZN (n_0_189_21), .A1 (n_0_189_6), .A2 (n_0_189_5), .A3 (n_0_189_4), .A4 (sps__n106));
INV_X1 i_0_189_12 (.ZN (n_0_189_20), .A (n_0_189_21));
NOR2_X1 i_0_189_11 (.ZN (n_0_189_19), .A1 (n_0_189_10), .A2 (n_0_189_34));
INV_X1 i_0_189_33 (.ZN (n_0_189_18), .A (sps__n36));
INV_X1 i_0_189_32 (.ZN (n_0_189_17), .A (sps__n7));
INV_X1 i_0_189_31 (.ZN (n_0_189_16), .A (sps__n13));
INV_X1 i_0_189_30 (.ZN (n_0_189_15), .A (sps__n49));
NAND4_X1 i_0_189_4 (.ZN (n_0_189_14), .A1 (n_0_189_18), .A2 (n_0_189_17), .A3 (n_0_189_16), .A4 (n_0_189_15));
INV_X1 i_0_189_3 (.ZN (n_0_189_13), .A (sps__n61));
INV_X1 i_0_189_2 (.ZN (n_0_189_12), .A (sps__n73));
INV_X1 i_0_189_1 (.ZN (n_0_189_11), .A (sps__n85));
NAND4_X1 i_0_189_0 (.ZN (n_0_189_10), .A1 (n_0_189_13), .A2 (n_0_189_12), .A3 (n_0_189_11), .A4 (sps__n1));
INV_X1 i_0_189_20 (.ZN (n_0_189_9), .A (sps__n119));
INV_X1 i_0_189_19 (.ZN (n_0_189_8), .A (sps__n113));
INV_X1 i_0_189_18 (.ZN (n_0_189_7), .A (sps__n97));
INV_X1 i_0_189_15 (.ZN (n_0_189_6), .A (sps__n69));
INV_X1 i_0_189_14 (.ZN (n_0_189_5), .A (sps__n21));
INV_X1 i_0_189_13 (.ZN (n_0_189_4), .A (sps__n79));
INV_X1 i_0_189_10 (.ZN (n_0_189_3), .A (sps__n56));
INV_X1 i_0_189_9 (.ZN (n_0_189_2), .A (sps__n27));
INV_X1 i_0_189_8 (.ZN (n_0_189_1), .A (sps__n41));
INV_X1 i_0_189_7 (.ZN (n_0_189_0), .A (sps__n93));
INV_X1 i_0_66_2 (.ZN (n_0_66_1), .A (sps__n62));
NAND2_X1 i_0_66_1 (.ZN (n_0_66_0), .A1 (n_0_66_1), .A2 (sps__n74));
INV_X2 i_0_66_0 (.ZN (n_0_5), .A (n_0_66_0));
INV_X1 i_0_49_39 (.ZN (n_0_49_38), .A (sps__n114));
INV_X1 i_0_49_38 (.ZN (n_0_49_37), .A (sps__n123));
INV_X1 i_0_49_37 (.ZN (n_0_49_36), .A (\mem[9][9] ));
NAND2_X1 i_0_49_36 (.ZN (n_0_49_35), .A1 (sps__n103), .A2 (n_0_49_36));
INV_X1 i_0_49_35 (.ZN (n_0_49_34), .A (sps__n103));
INV_X1 i_0_49_34 (.ZN (n_0_49_33), .A (\mem[1][9] ));
NAND2_X1 i_0_49_33 (.ZN (n_0_49_32), .A1 (n_0_49_34), .A2 (n_0_49_33));
NAND3_X1 i_0_49_32 (.ZN (n_0_49_31), .A1 (n_0_49_32), .A2 (n_0_49_37), .A3 (n_0_49_35));
NAND3_X1 i_0_49_31 (.ZN (n_0_49_30), .A1 (n_0_49_34), .A2 (sps__n123), .A3 (\mem[5][9] ));
NAND2_X1 i_0_49_30 (.ZN (n_0_49_29), .A1 (n_0_49_31), .A2 (n_0_49_30));
NAND2_X1 i_0_49_29 (.ZN (n_0_49_28), .A1 (n_0_49_29), .A2 (n_0_49_38));
NAND2_X1 i_0_49_28 (.ZN (n_0_49_27), .A1 (n_0_49_34), .A2 (sps__n114));
INV_X1 i_0_49_27 (.ZN (n_0_49_26), .A (n_0_49_27));
NAND2_X1 i_0_49_26 (.ZN (n_0_49_25), .A1 (n_0_49_4), .A2 (n_0_49_26));
NAND2_X1 i_0_49_25 (.ZN (n_0_49_24), .A1 (n_0_49_28), .A2 (n_0_49_25));
NOR2_X1 i_0_49_24 (.ZN (n_0_49_23), .A1 (n_0_49_1), .A2 (n_0_49_5));
NAND2_X1 i_0_49_23 (.ZN (n_0_49_22), .A1 (n_0_49_24), .A2 (n_0_49_23));
NAND2_X1 i_0_49_22 (.ZN (n_0_49_21), .A1 (sps__n103), .A2 (\mem[8][9] ));
NAND2_X1 i_0_49_21 (.ZN (n_0_49_20), .A1 (n_0_49_34), .A2 (\mem[0][9] ));
NAND3_X1 i_0_49_20 (.ZN (n_0_49_19), .A1 (n_0_49_20), .A2 (n_0_49_37), .A3 (n_0_49_21));
INV_X1 i_0_49_19 (.ZN (n_0_49_18), .A (\mem[4][9] ));
OAI21_X1 i_0_49_18 (.ZN (n_0_49_17), .A (sps__n123), .B1 (sps__n103), .B2 (n_0_49_18));
NAND3_X1 i_0_49_17 (.ZN (n_0_49_16), .A1 (n_0_49_19), .A2 (n_0_49_38), .A3 (n_0_49_17));
NAND2_X1 i_0_49_16 (.ZN (n_0_49_15), .A1 (sps__n103), .A2 (\mem[10][9] ));
NAND2_X1 i_0_49_15 (.ZN (n_0_49_14), .A1 (n_0_49_34), .A2 (\mem[2][9] ));
NAND3_X1 i_0_49_14 (.ZN (n_0_49_13), .A1 (n_0_49_14), .A2 (n_0_49_37), .A3 (n_0_49_15));
INV_X1 i_0_49_13 (.ZN (n_0_49_12), .A (\mem[6][9] ));
OAI21_X1 i_0_49_12 (.ZN (n_0_49_11), .A (sps__n123), .B1 (sps__n103), .B2 (n_0_49_12));
NAND3_X1 i_0_49_11 (.ZN (n_0_49_10), .A1 (n_0_49_13), .A2 (sps__n114), .A3 (n_0_49_11));
NAND2_X1 i_0_49_10 (.ZN (n_0_49_9), .A1 (n_0_49_16), .A2 (n_0_49_10));
NOR2_X1 i_0_49_9 (.ZN (n_0_49_8), .A1 (n_0_49_1), .A2 (sps__n98));
NAND2_X1 i_0_49_8 (.ZN (n_0_49_7), .A1 (n_0_49_9), .A2 (n_0_49_8));
NAND2_X1 i_0_49_7 (.ZN (n_0_49_6), .A1 (n_0_49_1), .A2 (dataout[9]));
NAND3_X1 i_0_49_6 (.ZN (n_0_4), .A1 (n_0_49_22), .A2 (n_0_49_7), .A3 (n_0_49_6));
INV_X1 i_0_49_5 (.ZN (n_0_49_5), .A (sps__n98));
NAND2_X1 i_0_49_4 (.ZN (n_0_49_4), .A1 (n_0_49_2), .A2 (n_0_49_3));
NAND2_X1 i_0_49_3 (.ZN (n_0_49_3), .A1 (sps__n123), .A2 (\mem[7][9] ));
NAND2_X1 i_0_49_2 (.ZN (n_0_49_2), .A1 (n_0_49_37), .A2 (\mem[3][9] ));
NAND2_X1 i_0_49_1 (.ZN (n_0_49_1), .A1 (n_0_49_0), .A2 (sps__n74));
INV_X1 i_0_49_0 (.ZN (n_0_49_0), .A (sps__n62));
NAND2_X1 i_0_7_39 (.ZN (n_0_7_38), .A1 (n_0_7_37), .A2 (\mem[9][0] ));
NAND2_X1 i_0_7_38 (.ZN (n_0_7_37), .A1 (n_0_7_0), .A2 (n_0_7_14));
NAND4_X1 i_0_7_37 (.ZN (n_0_7_36), .A1 (n_0_7_30), .A2 (n_0_7_32), .A3 (n_0_7_34), .A4 (n_0_7_35));
NOR2_X1 i_0_7_36 (.ZN (n_0_7_35), .A1 (sps__n112), .A2 (sps__n121));
INV_X1 i_0_7_35 (.ZN (n_0_7_34), .A (n_0_7_33));
NAND3_X1 i_0_7_34 (.ZN (n_0_7_33), .A1 (n_0_7_23), .A2 (sps__n97), .A3 (sps__n106));
INV_X1 i_0_7_33 (.ZN (n_0_7_32), .A (n_0_7_31));
NAND3_X1 i_0_7_28 (.ZN (n_0_7_31), .A1 (n_0_7_22), .A2 (n_0_7_21), .A3 (n_0_7_20));
INV_X1 i_0_7_27 (.ZN (n_0_7_30), .A (n_0_7_29));
NAND3_X1 i_0_7_23 (.ZN (n_0_7_29), .A1 (n_0_7_26), .A2 (n_0_7_25), .A3 (n_0_7_24));
INV_X1 i_0_7_22 (.ZN (n_0_7_28), .A (sps__n112));
INV_X1 i_0_7_16 (.ZN (n_0_7_27), .A (sps__n121));
INV_X1 i_0_7_15 (.ZN (n_0_7_26), .A (sps__n93));
INV_X1 i_0_7_14 (.ZN (n_0_7_25), .A (sps__n44));
INV_X1 i_0_7_13 (.ZN (n_0_7_24), .A (sps__n27));
INV_X1 i_0_7_12 (.ZN (n_0_7_23), .A (sps__n57));
INV_X1 i_0_7_11 (.ZN (n_0_7_22), .A (sps__n80));
INV_X1 i_0_7_10 (.ZN (n_0_7_21), .A (sps__n21));
INV_X1 i_0_7_21 (.ZN (n_0_7_20), .A (sps__n67));
NAND3_X1 i_0_7_8 (.ZN (n_0_7_19), .A1 (n_0_7_27), .A2 (n_0_7_28), .A3 (sps__n97));
NAND4_X1 i_0_7_20 (.ZN (n_0_7_18), .A1 (n_0_7_23), .A2 (n_0_7_24), .A3 (n_0_7_25), .A4 (n_0_7_26));
NAND4_X1 i_0_7_19 (.ZN (n_0_7_17), .A1 (n_0_7_20), .A2 (n_0_7_21), .A3 (n_0_7_22), .A4 (sps__n106));
INV_X1 i_0_7_2 (.ZN (n_0_7_16), .A (n_0_7_19));
NOR2_X1 i_0_7_18 (.ZN (n_0_7_15), .A1 (n_0_7_5), .A2 (n_0_7_18));
INV_X1 i_0_7_17 (.ZN (n_0_7_14), .A (n_0_7_5));
NAND2_X1 i_0_7_9 (.ZN (n_0_7_13), .A1 (n_0_7_36), .A2 (\mem[9][0] ));
NAND3_X1 i_0_7_7 (.ZN (n_0_7_12), .A1 (n_0_7_11), .A2 (n_0_7_15), .A3 (n_0_7_0));
NOR2_X1 i_0_7_6 (.ZN (n_0_7_11), .A1 (n_0_7_17), .A2 (n_0_7_10));
NAND2_X1 i_0_7_5 (.ZN (n_0_7_10), .A1 (n_0_7_16), .A2 (data[0]));
NAND3_X1 i_0_7_4 (.ZN (n_0_187), .A1 (n_0_7_12), .A2 (n_0_7_13), .A3 (n_0_7_38));
INV_X1 i_0_7_32 (.ZN (n_0_7_9), .A (sps__n35));
INV_X1 i_0_7_31 (.ZN (n_0_7_8), .A (sps__n8));
INV_X1 i_0_7_30 (.ZN (n_0_7_7), .A (sps__n13));
INV_X1 i_0_7_29 (.ZN (n_0_7_6), .A (sps__n49));
NAND4_X1 i_0_7_3 (.ZN (n_0_7_5), .A1 (n_0_7_9), .A2 (n_0_7_8), .A3 (n_0_7_7), .A4 (n_0_7_6));
INV_X1 i_0_7_26 (.ZN (n_0_7_4), .A (sps__n61));
INV_X1 i_0_7_25 (.ZN (n_0_7_3), .A (sps__n73));
INV_X1 i_0_7_24 (.ZN (n_0_7_2), .A (sps__n85));
NAND4_X1 i_0_7_1 (.ZN (n_0_7_1), .A1 (n_0_7_4), .A2 (n_0_7_3), .A3 (n_0_7_2), .A4 (sps__n1));
INV_X1 i_0_7_0 (.ZN (n_0_7_0), .A (n_0_7_1));
NOR2_X1 i_0_32_34 (.ZN (n_0_32_33), .A1 (n_0_32_19), .A2 (n_0_32_0));
INV_X1 i_0_32_33 (.ZN (n_0_32_32), .A (n_0_32_0));
INV_X1 i_0_32_28 (.ZN (n_0_32_31), .A (n_0_32_19));
NAND2_X1 i_0_32_27 (.ZN (n_0_32_30), .A1 (n_0_32_29), .A2 (\mem[10][0] ));
NAND3_X1 i_0_32_23 (.ZN (n_0_32_29), .A1 (n_0_32_5), .A2 (n_0_32_32), .A3 (n_0_32_10));
NAND3_X1 i_0_32_22 (.ZN (n_0_32_28), .A1 (n_0_32_27), .A2 (n_0_32_33), .A3 (n_0_32_14));
NOR2_X1 i_0_32_21 (.ZN (n_0_32_27), .A1 (n_0_32_6), .A2 (n_0_32_26));
NAND2_X1 i_0_32_20 (.ZN (n_0_32_26), .A1 (n_0_32_10), .A2 (data[0]));
NAND2_X1 i_0_32_19 (.ZN (n_0_32_25), .A1 (n_0_32_31), .A2 (n_0_32_14));
NAND3_X1 i_0_32_18 (.ZN (n_0_185), .A1 (n_0_32_28), .A2 (n_0_32_30), .A3 (n_0_32_24));
NAND2_X1 i_0_32_17 (.ZN (n_0_32_24), .A1 (n_0_32_25), .A2 (\mem[10][0] ));
INV_X1 i_0_32_32 (.ZN (n_0_32_23), .A (sps__n36));
INV_X1 i_0_32_31 (.ZN (n_0_32_22), .A (sps__n7));
INV_X1 i_0_32_30 (.ZN (n_0_32_21), .A (sps__n13));
INV_X1 i_0_32_29 (.ZN (n_0_32_20), .A (sps__n49));
NAND4_X1 i_0_32_3 (.ZN (n_0_32_19), .A1 (n_0_32_23), .A2 (n_0_32_22), .A3 (n_0_32_21), .A4 (n_0_32_20));
INV_X1 i_0_32_26 (.ZN (n_0_32_18), .A (sps__n61));
INV_X1 i_0_32_25 (.ZN (n_0_32_17), .A (sps__n73));
INV_X1 i_0_32_24 (.ZN (n_0_32_16), .A (sps__n85));
NAND4_X1 i_0_32_6 (.ZN (n_0_32_15), .A1 (n_0_32_18), .A2 (n_0_32_17), .A3 (n_0_32_16), .A4 (sps__n1));
INV_X1 i_0_32_16 (.ZN (n_0_32_14), .A (n_0_32_15));
INV_X1 i_0_32_15 (.ZN (n_0_32_13), .A (sps__n119));
INV_X1 i_0_32_14 (.ZN (n_0_32_12), .A (sps__n97));
NAND3_X1 i_0_32_13 (.ZN (n_0_32_11), .A1 (n_0_32_13), .A2 (n_0_32_12), .A3 (sps__n113));
INV_X1 i_0_32_12 (.ZN (n_0_32_10), .A (n_0_32_11));
INV_X1 i_0_32_11 (.ZN (n_0_32_9), .A (sps__n69));
INV_X1 i_0_32_10 (.ZN (n_0_32_8), .A (sps__n21));
INV_X1 i_0_32_9 (.ZN (n_0_32_7), .A (sps__n79));
NAND4_X1 i_0_32_8 (.ZN (n_0_32_6), .A1 (n_0_32_9), .A2 (n_0_32_8), .A3 (n_0_32_7), .A4 (sps__n103));
INV_X1 i_0_32_7 (.ZN (n_0_32_5), .A (n_0_32_6));
INV_X1 i_0_32_5 (.ZN (n_0_32_4), .A (sps__n56));
INV_X1 i_0_32_4 (.ZN (n_0_32_3), .A (sps__n27));
INV_X1 i_0_32_2 (.ZN (n_0_32_2), .A (sps__n41));
INV_X1 i_0_32_1 (.ZN (n_0_32_1), .A (sps__n93));
NAND4_X1 i_0_32_0 (.ZN (n_0_32_0), .A1 (n_0_32_4), .A2 (n_0_32_3), .A3 (n_0_32_2), .A4 (n_0_32_1));
INV_X1 i_0_190_39 (.ZN (n_0_190_38), .A (sps__n112));
INV_X1 i_0_190_38 (.ZN (n_0_190_37), .A (sps__n122));
INV_X1 i_0_190_37 (.ZN (n_0_190_36), .A (\mem[9][10] ));
NAND2_X1 i_0_190_36 (.ZN (n_0_190_35), .A1 (sps__n105), .A2 (n_0_190_36));
INV_X1 i_0_190_35 (.ZN (n_0_190_34), .A (sps__n105));
INV_X1 i_0_190_34 (.ZN (n_0_190_33), .A (\mem[1][10] ));
NAND2_X1 i_0_190_33 (.ZN (n_0_190_32), .A1 (n_0_190_34), .A2 (n_0_190_33));
NAND3_X1 i_0_190_32 (.ZN (n_0_190_31), .A1 (n_0_190_32), .A2 (n_0_190_37), .A3 (n_0_190_35));
NAND3_X1 i_0_190_31 (.ZN (n_0_190_30), .A1 (n_0_190_34), .A2 (sps__n122), .A3 (\mem[5][10] ));
NAND2_X1 i_0_190_30 (.ZN (n_0_190_29), .A1 (n_0_190_31), .A2 (n_0_190_30));
NAND2_X1 i_0_190_29 (.ZN (n_0_190_28), .A1 (n_0_190_29), .A2 (n_0_190_38));
NAND2_X1 i_0_190_28 (.ZN (n_0_190_27), .A1 (n_0_190_34), .A2 (sps__n112));
INV_X1 i_0_190_27 (.ZN (n_0_190_26), .A (n_0_190_27));
NAND2_X1 i_0_190_26 (.ZN (n_0_190_25), .A1 (n_0_190_4), .A2 (n_0_190_26));
NAND2_X1 i_0_190_25 (.ZN (n_0_190_24), .A1 (n_0_190_28), .A2 (n_0_190_25));
NOR2_X1 i_0_190_24 (.ZN (n_0_190_23), .A1 (n_0_190_1), .A2 (n_0_190_5));
NAND2_X1 i_0_190_23 (.ZN (n_0_190_22), .A1 (n_0_190_24), .A2 (n_0_190_23));
NAND2_X1 i_0_190_22 (.ZN (n_0_190_21), .A1 (sps__n105), .A2 (\mem[8][10] ));
NAND2_X1 i_0_190_21 (.ZN (n_0_190_20), .A1 (n_0_190_34), .A2 (\mem[0][10] ));
NAND3_X1 i_0_190_20 (.ZN (n_0_190_19), .A1 (n_0_190_20), .A2 (n_0_190_37), .A3 (n_0_190_21));
INV_X1 i_0_190_19 (.ZN (n_0_190_18), .A (\mem[4][10] ));
OAI21_X1 i_0_190_18 (.ZN (n_0_190_17), .A (sps__n122), .B1 (sps__n105), .B2 (n_0_190_18));
NAND3_X1 i_0_190_17 (.ZN (n_0_190_16), .A1 (n_0_190_19), .A2 (n_0_190_38), .A3 (n_0_190_17));
NAND2_X1 i_0_190_16 (.ZN (n_0_190_15), .A1 (sps__n105), .A2 (\mem[10][10] ));
NAND2_X1 i_0_190_15 (.ZN (n_0_190_14), .A1 (n_0_190_34), .A2 (\mem[2][10] ));
NAND3_X1 i_0_190_14 (.ZN (n_0_190_13), .A1 (n_0_190_14), .A2 (n_0_190_37), .A3 (n_0_190_15));
INV_X1 i_0_190_13 (.ZN (n_0_190_12), .A (\mem[6][10] ));
OAI21_X1 i_0_190_12 (.ZN (n_0_190_11), .A (sps__n122), .B1 (sps__n105), .B2 (n_0_190_12));
NAND3_X1 i_0_190_11 (.ZN (n_0_190_10), .A1 (n_0_190_13), .A2 (sps__n112), .A3 (n_0_190_11));
NAND2_X1 i_0_190_10 (.ZN (n_0_190_9), .A1 (n_0_190_16), .A2 (n_0_190_10));
NOR2_X1 i_0_190_9 (.ZN (n_0_190_8), .A1 (n_0_190_1), .A2 (sps__n99));
NAND2_X1 i_0_190_8 (.ZN (n_0_190_7), .A1 (n_0_190_9), .A2 (n_0_190_8));
NAND2_X1 i_0_190_7 (.ZN (n_0_190_6), .A1 (n_0_190_1), .A2 (dataout[10]));
NAND3_X1 i_0_190_6 (.ZN (n_0_151), .A1 (n_0_190_22), .A2 (n_0_190_7), .A3 (n_0_190_6));
INV_X1 i_0_190_5 (.ZN (n_0_190_5), .A (sps__n99));
NAND2_X1 i_0_190_4 (.ZN (n_0_190_4), .A1 (n_0_190_2), .A2 (n_0_190_3));
NAND2_X1 i_0_190_3 (.ZN (n_0_190_3), .A1 (sps__n122), .A2 (\mem[7][10] ));
NAND2_X1 i_0_190_2 (.ZN (n_0_190_2), .A1 (n_0_190_37), .A2 (\mem[3][10] ));
NAND2_X1 i_0_190_1 (.ZN (n_0_190_1), .A1 (n_0_190_0), .A2 (sps__n75));
INV_X1 i_0_190_0 (.ZN (n_0_190_0), .A (sps__n62));
NOR2_X1 i_0_6_34 (.ZN (n_0_6_33), .A1 (n_0_6_19), .A2 (n_0_6_0));
INV_X1 i_0_6_33 (.ZN (n_0_6_32), .A (n_0_6_0));
INV_X1 i_0_6_28 (.ZN (n_0_6_31), .A (n_0_6_19));
NAND2_X1 i_0_6_27 (.ZN (n_0_6_30), .A1 (n_0_6_29), .A2 (\mem[9][1] ));
NAND3_X1 i_0_6_23 (.ZN (n_0_6_29), .A1 (n_0_6_5), .A2 (n_0_6_32), .A3 (n_0_6_10));
NAND3_X1 i_0_6_22 (.ZN (n_0_6_28), .A1 (n_0_6_27), .A2 (n_0_6_33), .A3 (n_0_6_14));
NOR2_X1 i_0_6_21 (.ZN (n_0_6_27), .A1 (n_0_6_6), .A2 (n_0_6_26));
NAND2_X1 i_0_6_20 (.ZN (n_0_6_26), .A1 (n_0_6_10), .A2 (data[1]));
NAND2_X1 i_0_6_19 (.ZN (n_0_6_25), .A1 (n_0_6_31), .A2 (n_0_6_14));
NAND3_X1 i_0_6_18 (.ZN (n_0_150), .A1 (n_0_6_28), .A2 (n_0_6_30), .A3 (n_0_6_24));
NAND2_X1 i_0_6_17 (.ZN (n_0_6_24), .A1 (n_0_6_25), .A2 (\mem[9][1] ));
INV_X1 i_0_6_32 (.ZN (n_0_6_23), .A (sps__n34));
INV_X1 i_0_6_31 (.ZN (n_0_6_22), .A (sps__n7));
INV_X1 i_0_6_30 (.ZN (n_0_6_21), .A (sps__n13));
INV_X1 i_0_6_29 (.ZN (n_0_6_20), .A (sps__n49));
NAND4_X1 i_0_6_3 (.ZN (n_0_6_19), .A1 (n_0_6_23), .A2 (n_0_6_22), .A3 (n_0_6_21), .A4 (n_0_6_20));
INV_X1 i_0_6_26 (.ZN (n_0_6_18), .A (sps__n61));
INV_X1 i_0_6_25 (.ZN (n_0_6_17), .A (sps__n73));
INV_X1 i_0_6_24 (.ZN (n_0_6_16), .A (sps__n85));
NAND4_X1 i_0_6_6 (.ZN (n_0_6_15), .A1 (n_0_6_18), .A2 (n_0_6_17), .A3 (n_0_6_16), .A4 (sps__n1));
INV_X1 i_0_6_16 (.ZN (n_0_6_14), .A (n_0_6_15));
INV_X1 i_0_6_15 (.ZN (n_0_6_13), .A (sps__n119));
INV_X1 i_0_6_14 (.ZN (n_0_6_12), .A (sps__n113));
NAND3_X1 i_0_6_13 (.ZN (n_0_6_11), .A1 (n_0_6_13), .A2 (n_0_6_12), .A3 (sps__n97));
INV_X1 i_0_6_12 (.ZN (n_0_6_10), .A (n_0_6_11));
INV_X1 i_0_6_11 (.ZN (n_0_6_9), .A (sps__n69));
INV_X1 i_0_6_10 (.ZN (n_0_6_8), .A (sps__n21));
INV_X1 i_0_6_9 (.ZN (n_0_6_7), .A (sps__n79));
NAND4_X1 i_0_6_8 (.ZN (n_0_6_6), .A1 (n_0_6_9), .A2 (n_0_6_8), .A3 (n_0_6_7), .A4 (sps__n103));
INV_X1 i_0_6_7 (.ZN (n_0_6_5), .A (n_0_6_6));
INV_X1 i_0_6_5 (.ZN (n_0_6_4), .A (sps__n56));
INV_X1 i_0_6_4 (.ZN (n_0_6_3), .A (sps__n27));
INV_X1 i_0_6_2 (.ZN (n_0_6_2), .A (sps__n41));
INV_X1 i_0_6_1 (.ZN (n_0_6_1), .A (sps__n93));
NAND4_X1 i_0_6_0 (.ZN (n_0_6_0), .A1 (n_0_6_4), .A2 (n_0_6_3), .A3 (n_0_6_2), .A4 (n_0_6_1));
NOR2_X1 i_0_48_34 (.ZN (n_0_48_33), .A1 (n_0_48_19), .A2 (n_0_48_0));
INV_X1 i_0_48_33 (.ZN (n_0_48_32), .A (n_0_48_0));
INV_X1 i_0_48_28 (.ZN (n_0_48_31), .A (n_0_48_19));
NAND2_X1 i_0_48_27 (.ZN (n_0_48_30), .A1 (n_0_48_29), .A2 (\mem[10][1] ));
NAND3_X1 i_0_48_23 (.ZN (n_0_48_29), .A1 (n_0_48_5), .A2 (n_0_48_32), .A3 (n_0_48_10));
NAND3_X1 i_0_48_22 (.ZN (n_0_48_28), .A1 (n_0_48_27), .A2 (n_0_48_33), .A3 (n_0_48_14));
NOR2_X1 i_0_48_21 (.ZN (n_0_48_27), .A1 (n_0_48_6), .A2 (n_0_48_26));
NAND2_X1 i_0_48_20 (.ZN (n_0_48_26), .A1 (n_0_48_10), .A2 (data[1]));
NAND2_X1 i_0_48_19 (.ZN (n_0_48_25), .A1 (n_0_48_31), .A2 (n_0_48_14));
NAND3_X1 i_0_48_18 (.ZN (n_0_117), .A1 (n_0_48_28), .A2 (n_0_48_30), .A3 (n_0_48_24));
NAND2_X1 i_0_48_17 (.ZN (n_0_48_24), .A1 (n_0_48_25), .A2 (\mem[10][1] ));
INV_X1 i_0_48_32 (.ZN (n_0_48_23), .A (sps__n34));
INV_X1 i_0_48_31 (.ZN (n_0_48_22), .A (sps__n7));
INV_X1 i_0_48_30 (.ZN (n_0_48_21), .A (sps__n13));
INV_X1 i_0_48_29 (.ZN (n_0_48_20), .A (sps__n49));
NAND4_X1 i_0_48_3 (.ZN (n_0_48_19), .A1 (n_0_48_23), .A2 (n_0_48_22), .A3 (n_0_48_21), .A4 (n_0_48_20));
INV_X1 i_0_48_26 (.ZN (n_0_48_18), .A (sps__n61));
INV_X1 i_0_48_25 (.ZN (n_0_48_17), .A (sps__n73));
INV_X1 i_0_48_24 (.ZN (n_0_48_16), .A (sps__n85));
NAND4_X1 i_0_48_6 (.ZN (n_0_48_15), .A1 (n_0_48_18), .A2 (n_0_48_17), .A3 (n_0_48_16), .A4 (sps__n1));
INV_X1 i_0_48_16 (.ZN (n_0_48_14), .A (n_0_48_15));
INV_X1 i_0_48_15 (.ZN (n_0_48_13), .A (sps__n119));
INV_X1 i_0_48_14 (.ZN (n_0_48_12), .A (sps__n97));
NAND3_X1 i_0_48_13 (.ZN (n_0_48_11), .A1 (n_0_48_13), .A2 (n_0_48_12), .A3 (sps__n113));
INV_X1 i_0_48_12 (.ZN (n_0_48_10), .A (n_0_48_11));
INV_X1 i_0_48_11 (.ZN (n_0_48_9), .A (sps__n69));
INV_X1 i_0_48_10 (.ZN (n_0_48_8), .A (sps__n21));
INV_X1 i_0_48_9 (.ZN (n_0_48_7), .A (sps__n79));
NAND4_X1 i_0_48_8 (.ZN (n_0_48_6), .A1 (n_0_48_9), .A2 (n_0_48_8), .A3 (n_0_48_7), .A4 (sps__n103));
INV_X1 i_0_48_7 (.ZN (n_0_48_5), .A (n_0_48_6));
INV_X1 i_0_48_5 (.ZN (n_0_48_4), .A (sps__n56));
INV_X1 i_0_48_4 (.ZN (n_0_48_3), .A (sps__n27));
INV_X1 i_0_48_2 (.ZN (n_0_48_2), .A (sps__n41));
INV_X1 i_0_48_1 (.ZN (n_0_48_1), .A (sps__n93));
NAND4_X1 i_0_48_0 (.ZN (n_0_48_0), .A1 (n_0_48_4), .A2 (n_0_48_3), .A3 (n_0_48_2), .A4 (n_0_48_1));
NOR2_X1 i_0_187_31 (.ZN (n_0_116), .A1 (n_0_187_29), .A2 (n_0_187_30));
NAND3_X1 i_0_187_30 (.ZN (n_0_187_30), .A1 (n_0_187_24), .A2 (n_0_187_18), .A3 (n_0_187_28));
NAND3_X1 i_0_187_29 (.ZN (n_0_187_29), .A1 (n_0_187_20), .A2 (n_0_187_26), .A3 (n_0_187_22));
INV_X1 i_0_187_28 (.ZN (n_0_187_28), .A (n_0_187_27));
NAND2_X1 i_0_187_27 (.ZN (n_0_187_27), .A1 (n_0_187_0), .A2 (n_0_187_4));
INV_X1 i_0_187_24 (.ZN (n_0_187_26), .A (n_0_187_25));
NAND3_X1 i_0_187_23 (.ZN (n_0_187_25), .A1 (n_0_187_1), .A2 (n_0_187_5), .A3 (n_0_187_3));
INV_X1 i_0_187_19 (.ZN (n_0_187_24), .A (n_0_187_23));
NAND3_X1 i_0_187_18 (.ZN (n_0_187_23), .A1 (n_0_187_2), .A2 (n_0_187_6), .A3 (n_0_187_7));
INV_X1 i_0_187_17 (.ZN (n_0_187_22), .A (n_0_187_21));
NAND3_X1 i_0_187_15 (.ZN (n_0_187_21), .A1 (n_0_187_13), .A2 (n_0_187_10), .A3 (n_0_187_11));
INV_X1 i_0_187_14 (.ZN (n_0_187_20), .A (n_0_187_19));
NAND3_X1 i_0_187_13 (.ZN (n_0_187_19), .A1 (n_0_187_8), .A2 (n_0_187_12), .A3 (n_0_187_9));
NOR2_X1 i_0_187_12 (.ZN (n_0_187_18), .A1 (n_0_187_16), .A2 (n_0_187_17));
NAND3_X1 i_0_187_10 (.ZN (n_0_187_17), .A1 (sps__n113), .A2 (address[0]), .A3 (sps__n1));
NAND2_X1 i_0_187_9 (.ZN (n_0_187_16), .A1 (n_0_187_14), .A2 (n_0_187_15));
INV_X1 i_0_187_8 (.ZN (n_0_187_15), .A (sps__n34));
INV_X1 i_0_187_6 (.ZN (n_0_187_14), .A (sps__n7));
INV_X1 i_0_187_26 (.ZN (n_0_187_13), .A (sps__n13));
INV_X1 i_0_187_25 (.ZN (n_0_187_12), .A (sps__n49));
INV_X1 i_0_187_22 (.ZN (n_0_187_11), .A (sps__n61));
INV_X1 i_0_187_21 (.ZN (n_0_187_10), .A (sps__n73));
INV_X1 i_0_187_20 (.ZN (n_0_187_9), .A (sps__n85));
INV_X1 i_0_187_16 (.ZN (n_0_187_8), .A (sps__n119));
INV_X1 i_0_187_4 (.ZN (n_0_187_7), .A (sps__n67));
INV_X1 i_0_187_3 (.ZN (n_0_187_6), .A (sps__n21));
INV_X1 i_0_187_11 (.ZN (n_0_187_5), .A (sps__n79));
INV_X1 i_0_187_2 (.ZN (n_0_187_4), .A (sps__n106));
INV_X1 i_0_187_7 (.ZN (n_0_187_3), .A (sps__n56));
INV_X1 i_0_187_1 (.ZN (n_0_187_2), .A (sps__n27));
INV_X1 i_0_187_5 (.ZN (n_0_187_1), .A (sps__n41));
INV_X1 i_0_187_0 (.ZN (n_0_187_0), .A (sps__n93));
NAND3_X1 i_0_31_31 (.ZN (n_0_31_30), .A1 (n_0_31_27), .A2 (n_0_31_28), .A3 (n_0_31_29));
NOR2_X1 i_0_31_30 (.ZN (n_0_31_29), .A1 (n_0_31_13), .A2 (n_0_31_23));
NOR2_X1 i_0_31_29 (.ZN (n_0_31_28), .A1 (n_0_31_22), .A2 (n_0_31_21));
NOR2_X1 i_0_31_28 (.ZN (n_0_31_27), .A1 (n_0_31_17), .A2 (n_0_31_20));
NOR2_X1 i_0_31_27 (.ZN (n_0_31_26), .A1 (n_0_31_17), .A2 (n_0_31_13));
NOR2_X1 i_0_31_26 (.ZN (n_0_31_25), .A1 (n_0_31_20), .A2 (n_0_31_21));
NOR2_X1 i_0_31_25 (.ZN (n_0_31_24), .A1 (n_0_31_22), .A2 (n_0_31_23));
NAND3_X1 i_0_31_24 (.ZN (n_0_31_23), .A1 (n_0_31_4), .A2 (n_0_31_2), .A3 (n_0_31_6));
NAND3_X1 i_0_31_23 (.ZN (n_0_31_22), .A1 (n_0_31_1), .A2 (n_0_31_3), .A3 (n_0_31_5));
NAND3_X1 i_0_31_22 (.ZN (n_0_31_21), .A1 (n_0_31_10), .A2 (n_0_31_8), .A3 (n_0_31_12));
NAND3_X1 i_0_31_21 (.ZN (n_0_31_20), .A1 (n_0_31_7), .A2 (n_0_31_9), .A3 (n_0_31_11));
NAND2_X1 i_0_31_20 (.ZN (n_0_31_19), .A1 (n_0_31_30), .A2 (\mem[3][1] ));
INV_X1 i_0_31_19 (.ZN (n_0_31_18), .A (sps__n119));
NAND4_X1 i_0_31_18 (.ZN (n_0_31_17), .A1 (n_0_31_18), .A2 (sps__n1), .A3 (sps__n113), .A4 (address[0]));
INV_X1 i_0_31_17 (.ZN (n_0_31_16), .A (sps__n21));
INV_X1 i_0_31_16 (.ZN (n_0_31_15), .A (sps__n79));
INV_X1 i_0_31_15 (.ZN (n_0_31_14), .A (sps__n106));
NAND3_X1 i_0_31_14 (.ZN (n_0_31_13), .A1 (n_0_31_16), .A2 (n_0_31_15), .A3 (n_0_31_14));
INV_X1 i_0_31_13 (.ZN (n_0_31_12), .A (sps__n61));
INV_X1 i_0_31_12 (.ZN (n_0_31_11), .A (sps__n73));
INV_X1 i_0_31_11 (.ZN (n_0_31_10), .A (sps__n7));
INV_X1 i_0_31_10 (.ZN (n_0_31_9), .A (sps__n13));
INV_X1 i_0_31_9 (.ZN (n_0_31_8), .A (sps__n85));
INV_X1 i_0_31_8 (.ZN (n_0_31_7), .A (sps__n34));
INV_X1 i_0_31_7 (.ZN (n_0_31_6), .A (sps__n93));
INV_X1 i_0_31_6 (.ZN (n_0_31_5), .A (sps__n69));
INV_X1 i_0_31_5 (.ZN (n_0_31_4), .A (sps__n27));
INV_X1 i_0_31_4 (.ZN (n_0_31_3), .A (sps__n41));
INV_X1 i_0_31_3 (.ZN (n_0_31_2), .A (sps__n49));
INV_X1 i_0_31_2 (.ZN (n_0_31_1), .A (sps__n56));
NAND4_X1 i_0_31_1 (.ZN (n_0_31_0), .A1 (n_0_31_26), .A2 (n_0_31_25), .A3 (n_0_31_24), .A4 (data[1]));
NAND2_X1 i_0_31_0 (.ZN (n_0_100), .A1 (n_0_31_19), .A2 (n_0_31_0));
NOR2_X1 i_0_150_31 (.ZN (n_0_99), .A1 (n_0_150_29), .A2 (n_0_150_30));
NAND3_X1 i_0_150_30 (.ZN (n_0_150_30), .A1 (n_0_150_24), .A2 (n_0_150_18), .A3 (n_0_150_28));
NAND3_X1 i_0_150_29 (.ZN (n_0_150_29), .A1 (n_0_150_20), .A2 (n_0_150_26), .A3 (n_0_150_22));
INV_X1 i_0_150_28 (.ZN (n_0_150_28), .A (n_0_150_27));
NAND2_X1 i_0_150_27 (.ZN (n_0_150_27), .A1 (n_0_150_0), .A2 (n_0_150_4));
INV_X1 i_0_150_24 (.ZN (n_0_150_26), .A (n_0_150_25));
NAND3_X1 i_0_150_23 (.ZN (n_0_150_25), .A1 (n_0_150_1), .A2 (n_0_150_5), .A3 (n_0_150_3));
INV_X1 i_0_150_19 (.ZN (n_0_150_24), .A (n_0_150_23));
NAND3_X1 i_0_150_18 (.ZN (n_0_150_23), .A1 (n_0_150_2), .A2 (n_0_150_6), .A3 (n_0_150_7));
INV_X1 i_0_150_17 (.ZN (n_0_150_22), .A (n_0_150_21));
NAND3_X1 i_0_150_15 (.ZN (n_0_150_21), .A1 (n_0_150_13), .A2 (n_0_150_10), .A3 (n_0_150_11));
INV_X1 i_0_150_14 (.ZN (n_0_150_20), .A (n_0_150_19));
NAND3_X1 i_0_150_13 (.ZN (n_0_150_19), .A1 (n_0_150_8), .A2 (n_0_150_12), .A3 (n_0_150_9));
NOR2_X1 i_0_150_12 (.ZN (n_0_150_18), .A1 (n_0_150_16), .A2 (n_0_150_17));
NAND3_X1 i_0_150_10 (.ZN (n_0_150_17), .A1 (sps__n121), .A2 (sps__n97), .A3 (sps__n1));
NAND2_X1 i_0_150_9 (.ZN (n_0_150_16), .A1 (n_0_150_14), .A2 (n_0_150_15));
INV_X1 i_0_150_8 (.ZN (n_0_150_15), .A (sps__n35));
INV_X1 i_0_150_6 (.ZN (n_0_150_14), .A (sps__n8));
INV_X1 i_0_150_26 (.ZN (n_0_150_13), .A (sps__n13));
INV_X1 i_0_150_25 (.ZN (n_0_150_12), .A (sps__n49));
INV_X1 i_0_150_22 (.ZN (n_0_150_11), .A (sps__n61));
INV_X1 i_0_150_21 (.ZN (n_0_150_10), .A (sps__n73));
INV_X1 i_0_150_20 (.ZN (n_0_150_9), .A (sps__n85));
INV_X1 i_0_150_16 (.ZN (n_0_150_8), .A (sps__n112));
INV_X1 i_0_150_4 (.ZN (n_0_150_7), .A (sps__n67));
INV_X1 i_0_150_3 (.ZN (n_0_150_6), .A (sps__n21));
INV_X1 i_0_150_11 (.ZN (n_0_150_5), .A (sps__n79));
INV_X1 i_0_150_2 (.ZN (n_0_150_4), .A (sps__n106));
INV_X1 i_0_150_7 (.ZN (n_0_150_3), .A (sps__n56));
INV_X1 i_0_150_1 (.ZN (n_0_150_2), .A (sps__n27));
INV_X1 i_0_150_5 (.ZN (n_0_150_1), .A (sps__n41));
INV_X1 i_0_150_0 (.ZN (n_0_150_0), .A (sps__n93));
NAND3_X1 i_0_149_31 (.ZN (n_0_149_30), .A1 (n_0_149_27), .A2 (n_0_149_28), .A3 (n_0_149_29));
NOR2_X1 i_0_149_30 (.ZN (n_0_149_29), .A1 (n_0_149_13), .A2 (n_0_149_23));
NOR2_X1 i_0_149_29 (.ZN (n_0_149_28), .A1 (n_0_149_22), .A2 (n_0_149_21));
NOR2_X1 i_0_149_28 (.ZN (n_0_149_27), .A1 (n_0_149_17), .A2 (n_0_149_20));
NOR2_X1 i_0_149_27 (.ZN (n_0_149_26), .A1 (n_0_149_17), .A2 (n_0_149_13));
NOR2_X1 i_0_149_26 (.ZN (n_0_149_25), .A1 (n_0_149_20), .A2 (n_0_149_21));
NOR2_X1 i_0_149_25 (.ZN (n_0_149_24), .A1 (n_0_149_22), .A2 (n_0_149_23));
NAND3_X1 i_0_149_24 (.ZN (n_0_149_23), .A1 (n_0_149_4), .A2 (n_0_149_2), .A3 (n_0_149_6));
NAND3_X1 i_0_149_23 (.ZN (n_0_149_22), .A1 (n_0_149_1), .A2 (n_0_149_3), .A3 (n_0_149_5));
NAND3_X1 i_0_149_22 (.ZN (n_0_149_21), .A1 (n_0_149_10), .A2 (n_0_149_8), .A3 (n_0_149_12));
NAND3_X1 i_0_149_21 (.ZN (n_0_149_20), .A1 (n_0_149_7), .A2 (n_0_149_9), .A3 (n_0_149_11));
NAND2_X1 i_0_149_20 (.ZN (n_0_149_19), .A1 (n_0_149_30), .A2 (\mem[5][1] ));
INV_X1 i_0_149_19 (.ZN (n_0_149_18), .A (sps__n113));
NAND4_X1 i_0_149_18 (.ZN (n_0_149_17), .A1 (n_0_149_18), .A2 (sps__n1), .A3 (sps__n119), .A4 (sps__n97));
INV_X1 i_0_149_17 (.ZN (n_0_149_16), .A (sps__n21));
INV_X1 i_0_149_16 (.ZN (n_0_149_15), .A (sps__n79));
INV_X1 i_0_149_15 (.ZN (n_0_149_14), .A (sps__n106));
NAND3_X1 i_0_149_14 (.ZN (n_0_149_13), .A1 (n_0_149_16), .A2 (n_0_149_15), .A3 (n_0_149_14));
INV_X1 i_0_149_13 (.ZN (n_0_149_12), .A (sps__n61));
INV_X1 i_0_149_12 (.ZN (n_0_149_11), .A (sps__n73));
INV_X1 i_0_149_11 (.ZN (n_0_149_10), .A (sps__n7));
INV_X1 i_0_149_10 (.ZN (n_0_149_9), .A (sps__n13));
INV_X1 i_0_149_9 (.ZN (n_0_149_8), .A (sps__n85));
INV_X1 i_0_149_8 (.ZN (n_0_149_7), .A (sps__n34));
INV_X1 i_0_149_7 (.ZN (n_0_149_6), .A (sps__n93));
INV_X1 i_0_149_6 (.ZN (n_0_149_5), .A (sps__n69));
INV_X1 i_0_149_5 (.ZN (n_0_149_4), .A (sps__n27));
INV_X1 i_0_149_4 (.ZN (n_0_149_3), .A (sps__n41));
INV_X1 i_0_149_3 (.ZN (n_0_149_2), .A (sps__n49));
INV_X1 i_0_149_2 (.ZN (n_0_149_1), .A (sps__n56));
NAND4_X1 i_0_149_1 (.ZN (n_0_149_0), .A1 (n_0_149_26), .A2 (n_0_149_25), .A3 (n_0_149_24), .A4 (data[1]));
NAND2_X1 i_0_149_0 (.ZN (n_0_66), .A1 (n_0_149_19), .A2 (n_0_149_0));
NOR2_X1 i_0_116_31 (.ZN (n_0_65), .A1 (n_0_116_29), .A2 (n_0_116_30));
NAND3_X1 i_0_116_30 (.ZN (n_0_116_30), .A1 (n_0_116_24), .A2 (n_0_116_18), .A3 (n_0_116_28));
NAND3_X1 i_0_116_29 (.ZN (n_0_116_29), .A1 (n_0_116_20), .A2 (n_0_116_26), .A3 (n_0_116_22));
INV_X1 i_0_116_28 (.ZN (n_0_116_28), .A (n_0_116_27));
NAND2_X1 i_0_116_27 (.ZN (n_0_116_27), .A1 (n_0_116_0), .A2 (n_0_116_4));
INV_X1 i_0_116_24 (.ZN (n_0_116_26), .A (n_0_116_25));
NAND3_X1 i_0_116_23 (.ZN (n_0_116_25), .A1 (n_0_116_1), .A2 (n_0_116_5), .A3 (n_0_116_3));
INV_X1 i_0_116_19 (.ZN (n_0_116_24), .A (n_0_116_23));
NAND3_X1 i_0_116_18 (.ZN (n_0_116_23), .A1 (n_0_116_2), .A2 (n_0_116_6), .A3 (n_0_116_7));
INV_X1 i_0_116_17 (.ZN (n_0_116_22), .A (n_0_116_21));
NAND3_X1 i_0_116_15 (.ZN (n_0_116_21), .A1 (n_0_116_13), .A2 (n_0_116_10), .A3 (n_0_116_11));
INV_X1 i_0_116_14 (.ZN (n_0_116_20), .A (n_0_116_19));
NAND3_X1 i_0_116_13 (.ZN (n_0_116_19), .A1 (n_0_116_8), .A2 (n_0_116_12), .A3 (n_0_116_9));
NOR2_X1 i_0_116_12 (.ZN (n_0_116_18), .A1 (n_0_116_16), .A2 (n_0_116_17));
NAND3_X1 i_0_116_10 (.ZN (n_0_116_17), .A1 (sps__n119), .A2 (sps__n113), .A3 (sps__n1));
NAND2_X1 i_0_116_9 (.ZN (n_0_116_16), .A1 (n_0_116_14), .A2 (n_0_116_15));
INV_X1 i_0_116_8 (.ZN (n_0_116_15), .A (sps__n34));
INV_X1 i_0_116_6 (.ZN (n_0_116_14), .A (sps__n7));
INV_X1 i_0_116_26 (.ZN (n_0_116_13), .A (sps__n13));
INV_X1 i_0_116_25 (.ZN (n_0_116_12), .A (sps__n49));
INV_X1 i_0_116_22 (.ZN (n_0_116_11), .A (sps__n61));
INV_X1 i_0_116_21 (.ZN (n_0_116_10), .A (sps__n73));
INV_X1 i_0_116_20 (.ZN (n_0_116_9), .A (sps__n85));
INV_X1 i_0_116_16 (.ZN (n_0_116_8), .A (sps__n97));
INV_X1 i_0_116_4 (.ZN (n_0_116_7), .A (sps__n67));
INV_X1 i_0_116_3 (.ZN (n_0_116_6), .A (sps__n21));
INV_X1 i_0_116_11 (.ZN (n_0_116_5), .A (sps__n79));
INV_X1 i_0_116_2 (.ZN (n_0_116_4), .A (sps__n106));
INV_X1 i_0_116_7 (.ZN (n_0_116_3), .A (sps__n56));
INV_X1 i_0_116_1 (.ZN (n_0_116_2), .A (sps__n27));
INV_X1 i_0_116_5 (.ZN (n_0_116_1), .A (sps__n41));
INV_X1 i_0_116_0 (.ZN (n_0_116_0), .A (sps__n93));
NAND3_X1 i_0_99_31 (.ZN (n_0_99_30), .A1 (n_0_99_27), .A2 (n_0_99_28), .A3 (n_0_99_29));
NOR2_X1 i_0_99_30 (.ZN (n_0_99_29), .A1 (n_0_99_13), .A2 (n_0_99_23));
NOR2_X1 i_0_99_29 (.ZN (n_0_99_28), .A1 (n_0_99_22), .A2 (n_0_99_21));
NOR2_X1 i_0_99_28 (.ZN (n_0_99_27), .A1 (n_0_99_17), .A2 (n_0_99_20));
NOR2_X1 i_0_99_27 (.ZN (n_0_99_26), .A1 (n_0_99_17), .A2 (n_0_99_13));
NOR2_X1 i_0_99_26 (.ZN (n_0_99_25), .A1 (n_0_99_20), .A2 (n_0_99_21));
NOR2_X1 i_0_99_25 (.ZN (n_0_99_24), .A1 (n_0_99_22), .A2 (n_0_99_23));
NAND3_X1 i_0_99_24 (.ZN (n_0_99_23), .A1 (n_0_99_4), .A2 (n_0_99_2), .A3 (n_0_99_6));
NAND3_X1 i_0_99_23 (.ZN (n_0_99_22), .A1 (n_0_99_1), .A2 (n_0_99_3), .A3 (n_0_99_5));
NAND3_X1 i_0_99_22 (.ZN (n_0_99_21), .A1 (n_0_99_10), .A2 (n_0_99_8), .A3 (n_0_99_12));
NAND3_X1 i_0_99_21 (.ZN (n_0_99_20), .A1 (n_0_99_7), .A2 (n_0_99_9), .A3 (n_0_99_11));
NAND2_X1 i_0_99_20 (.ZN (n_0_99_19), .A1 (n_0_99_30), .A2 (\mem[6][1] ));
INV_X1 i_0_99_19 (.ZN (n_0_99_18), .A (sps__n97));
NAND4_X1 i_0_99_18 (.ZN (n_0_99_17), .A1 (n_0_99_18), .A2 (sps__n1), .A3 (sps__n119), .A4 (sps__n113));
INV_X1 i_0_99_17 (.ZN (n_0_99_16), .A (sps__n21));
INV_X1 i_0_99_16 (.ZN (n_0_99_15), .A (sps__n79));
INV_X1 i_0_99_15 (.ZN (n_0_99_14), .A (sps__n106));
NAND3_X1 i_0_99_14 (.ZN (n_0_99_13), .A1 (n_0_99_16), .A2 (n_0_99_15), .A3 (n_0_99_14));
INV_X1 i_0_99_13 (.ZN (n_0_99_12), .A (sps__n61));
INV_X1 i_0_99_12 (.ZN (n_0_99_11), .A (sps__n73));
INV_X1 i_0_99_11 (.ZN (n_0_99_10), .A (sps__n7));
INV_X1 i_0_99_10 (.ZN (n_0_99_9), .A (sps__n13));
INV_X1 i_0_99_9 (.ZN (n_0_99_8), .A (sps__n85));
INV_X1 i_0_99_8 (.ZN (n_0_99_7), .A (sps__n34));
INV_X1 i_0_99_7 (.ZN (n_0_99_6), .A (sps__n93));
INV_X1 i_0_99_6 (.ZN (n_0_99_5), .A (sps__n69));
INV_X1 i_0_99_5 (.ZN (n_0_99_4), .A (sps__n27));
INV_X1 i_0_99_4 (.ZN (n_0_99_3), .A (sps__n41));
INV_X1 i_0_99_3 (.ZN (n_0_99_2), .A (sps__n49));
INV_X1 i_0_99_2 (.ZN (n_0_99_1), .A (sps__n56));
NAND4_X1 i_0_99_1 (.ZN (n_0_99_0), .A1 (n_0_99_26), .A2 (n_0_99_25), .A3 (n_0_99_24), .A4 (data[1]));
NAND2_X1 i_0_99_0 (.ZN (n_0_49), .A1 (n_0_99_19), .A2 (n_0_99_0));
DFF_X2 \temp_reg[9]  (.Q (dataout[9]), .CK (n_0_32), .D (n_0_4));
DFF_X2 \temp_reg[10]  (.Q (dataout[10]), .CK (n_0_32), .D (n_0_151));
DFF_X2 \mem_reg[3][0]  (.Q (\mem[3][0] ), .CK (n_0_32), .D (n_0_14));
DFF_X2 \mem_reg[3][1]  (.Q (\mem[3][1] ), .CK (n_0_32), .D (n_0_100));
DFF_X2 \mem_reg[5][0]  (.Q (\mem[5][0] ), .CK (n_0_32), .D (n_0_12));
DFF_X2 \mem_reg[5][1]  (.Q (\mem[5][1] ), .CK (n_0_32), .D (n_0_66));
DFF_X2 \mem_reg[6][0]  (.Q (\mem[6][0] ), .CK (n_0_32), .D (n_0_10));
DFF_X2 \mem_reg[6][1]  (.Q (\mem[6][1] ), .CK (n_0_32), .D (n_0_49));
DFF_X2 \temp_reg[5]  (.Q (dataout[5]), .CK (n_0_32), .D (n_0_16));
DFF_X2 \temp_reg[6]  (.Q (dataout[6]), .CK (n_0_32), .D (n_0_15));
NAND3_X1 i_0_193_31 (.ZN (n_0_193_30), .A1 (n_0_193_27), .A2 (n_0_193_28), .A3 (n_0_193_29));
NOR2_X1 i_0_193_30 (.ZN (n_0_193_29), .A1 (n_0_193_13), .A2 (n_0_193_23));
NOR2_X1 i_0_193_29 (.ZN (n_0_193_28), .A1 (n_0_193_22), .A2 (n_0_193_21));
NOR2_X1 i_0_193_28 (.ZN (n_0_193_27), .A1 (n_0_193_17), .A2 (n_0_193_20));
NOR2_X1 i_0_193_27 (.ZN (n_0_193_26), .A1 (n_0_193_17), .A2 (n_0_193_13));
NOR2_X1 i_0_193_26 (.ZN (n_0_193_25), .A1 (n_0_193_20), .A2 (n_0_193_21));
NOR2_X1 i_0_193_25 (.ZN (n_0_193_24), .A1 (n_0_193_22), .A2 (n_0_193_23));
NAND3_X1 i_0_193_24 (.ZN (n_0_193_23), .A1 (n_0_193_4), .A2 (n_0_193_2), .A3 (n_0_193_6));
NAND3_X1 i_0_193_23 (.ZN (n_0_193_22), .A1 (n_0_193_1), .A2 (n_0_193_3), .A3 (n_0_193_5));
NAND3_X1 i_0_193_22 (.ZN (n_0_193_21), .A1 (n_0_193_10), .A2 (n_0_193_8), .A3 (n_0_193_12));
NAND3_X1 i_0_193_21 (.ZN (n_0_193_20), .A1 (n_0_193_7), .A2 (n_0_193_9), .A3 (n_0_193_11));
NAND2_X1 i_0_193_20 (.ZN (n_0_193_19), .A1 (n_0_193_30), .A2 (\mem[3][2] ));
INV_X1 i_0_193_19 (.ZN (n_0_193_18), .A (sps__n121));
NAND4_X1 i_0_193_18 (.ZN (n_0_193_17), .A1 (n_0_193_18), .A2 (sps__n1), .A3 (sps__n112), .A4 (sps__n97));
INV_X1 i_0_193_17 (.ZN (n_0_193_16), .A (sps__n21));
INV_X1 i_0_193_16 (.ZN (n_0_193_15), .A (sps__n80));
INV_X1 i_0_193_15 (.ZN (n_0_193_14), .A (sps__n106));
NAND3_X1 i_0_193_14 (.ZN (n_0_193_13), .A1 (n_0_193_16), .A2 (n_0_193_15), .A3 (n_0_193_14));
INV_X1 i_0_193_13 (.ZN (n_0_193_12), .A (sps__n63));
INV_X1 i_0_193_12 (.ZN (n_0_193_11), .A (sps__n75));
INV_X1 i_0_193_11 (.ZN (n_0_193_10), .A (sps__n8));
INV_X1 i_0_193_10 (.ZN (n_0_193_9), .A (sps__n13));
INV_X1 i_0_193_9 (.ZN (n_0_193_8), .A (sps__n87));
INV_X1 i_0_193_8 (.ZN (n_0_193_7), .A (sps__n35));
INV_X1 i_0_193_7 (.ZN (n_0_193_6), .A (sps__n93));
INV_X1 i_0_193_6 (.ZN (n_0_193_5), .A (sps__n67));
INV_X1 i_0_193_5 (.ZN (n_0_193_4), .A (sps__n27));
INV_X1 i_0_193_4 (.ZN (n_0_193_3), .A (sps__n44));
INV_X1 i_0_193_3 (.ZN (n_0_193_2), .A (sps__n50));
INV_X1 i_0_193_2 (.ZN (n_0_193_1), .A (sps__n57));
NAND4_X1 i_0_193_1 (.ZN (n_0_193_0), .A1 (n_0_193_26), .A2 (n_0_193_25), .A3 (n_0_193_24), .A4 (data[2]));
NAND2_X1 i_0_193_0 (.ZN (n_0_3), .A1 (n_0_193_19), .A2 (n_0_193_0));
NAND3_X1 i_0_134_31 (.ZN (n_0_134_30), .A1 (n_0_134_27), .A2 (n_0_134_28), .A3 (n_0_134_29));
NOR2_X1 i_0_134_30 (.ZN (n_0_134_29), .A1 (n_0_134_13), .A2 (n_0_134_23));
NOR2_X1 i_0_134_29 (.ZN (n_0_134_28), .A1 (n_0_134_22), .A2 (n_0_134_21));
NOR2_X1 i_0_134_28 (.ZN (n_0_134_27), .A1 (n_0_134_17), .A2 (n_0_134_20));
NOR2_X1 i_0_134_27 (.ZN (n_0_134_26), .A1 (n_0_134_17), .A2 (n_0_134_13));
NOR2_X1 i_0_134_26 (.ZN (n_0_134_25), .A1 (n_0_134_20), .A2 (n_0_134_21));
NOR2_X1 i_0_134_25 (.ZN (n_0_134_24), .A1 (n_0_134_22), .A2 (n_0_134_23));
NAND3_X1 i_0_134_24 (.ZN (n_0_134_23), .A1 (n_0_134_4), .A2 (n_0_134_2), .A3 (n_0_134_6));
NAND3_X1 i_0_134_23 (.ZN (n_0_134_22), .A1 (n_0_134_1), .A2 (n_0_134_3), .A3 (n_0_134_5));
NAND3_X1 i_0_134_22 (.ZN (n_0_134_21), .A1 (n_0_134_10), .A2 (n_0_134_8), .A3 (n_0_134_12));
NAND3_X1 i_0_134_21 (.ZN (n_0_134_20), .A1 (n_0_134_7), .A2 (n_0_134_9), .A3 (n_0_134_11));
NAND2_X1 i_0_134_20 (.ZN (n_0_134_19), .A1 (n_0_134_30), .A2 (\mem[5][2] ));
INV_X1 i_0_134_19 (.ZN (n_0_134_18), .A (sps__n112));
NAND4_X1 i_0_134_18 (.ZN (n_0_134_17), .A1 (n_0_134_18), .A2 (sps__n3), .A3 (sps__n121), .A4 (sps__n99));
INV_X1 i_0_134_17 (.ZN (n_0_134_16), .A (sps__n21));
INV_X1 i_0_134_16 (.ZN (n_0_134_15), .A (sps__n80));
INV_X1 i_0_134_15 (.ZN (n_0_134_14), .A (sps__n103));
NAND3_X1 i_0_134_14 (.ZN (n_0_134_13), .A1 (n_0_134_16), .A2 (n_0_134_15), .A3 (n_0_134_14));
INV_X1 i_0_134_13 (.ZN (n_0_134_12), .A (sps__n63));
INV_X1 i_0_134_12 (.ZN (n_0_134_11), .A (sps__n74));
INV_X1 i_0_134_11 (.ZN (n_0_134_10), .A (sps__n8));
INV_X1 i_0_134_10 (.ZN (n_0_134_9), .A (sps__n13));
INV_X1 i_0_134_9 (.ZN (n_0_134_8), .A (sps__n87));
INV_X1 i_0_134_8 (.ZN (n_0_134_7), .A (sps__n35));
INV_X1 i_0_134_7 (.ZN (n_0_134_6), .A (sps__n93));
INV_X1 i_0_134_6 (.ZN (n_0_134_5), .A (sps__n67));
INV_X1 i_0_134_5 (.ZN (n_0_134_4), .A (sps__n27));
INV_X1 i_0_134_4 (.ZN (n_0_134_3), .A (sps__n44));
INV_X1 i_0_134_3 (.ZN (n_0_134_2), .A (sps__n49));
INV_X1 i_0_134_2 (.ZN (n_0_134_1), .A (sps__n57));
NAND4_X1 i_0_134_1 (.ZN (n_0_134_0), .A1 (n_0_134_26), .A2 (n_0_134_25), .A3 (n_0_134_24), .A4 (data[2]));
NAND2_X1 i_0_134_0 (.ZN (n_0_2), .A1 (n_0_134_19), .A2 (n_0_134_0));
NAND3_X1 i_0_115_31 (.ZN (n_0_115_30), .A1 (n_0_115_27), .A2 (n_0_115_28), .A3 (n_0_115_29));
NOR2_X1 i_0_115_30 (.ZN (n_0_115_29), .A1 (n_0_115_13), .A2 (n_0_115_23));
NOR2_X1 i_0_115_29 (.ZN (n_0_115_28), .A1 (n_0_115_22), .A2 (n_0_115_21));
NOR2_X1 i_0_115_28 (.ZN (n_0_115_27), .A1 (n_0_115_17), .A2 (n_0_115_20));
NOR2_X1 i_0_115_27 (.ZN (n_0_115_26), .A1 (n_0_115_17), .A2 (n_0_115_13));
NOR2_X1 i_0_115_26 (.ZN (n_0_115_25), .A1 (n_0_115_20), .A2 (n_0_115_21));
NOR2_X1 i_0_115_25 (.ZN (n_0_115_24), .A1 (n_0_115_22), .A2 (n_0_115_23));
NAND3_X1 i_0_115_24 (.ZN (n_0_115_23), .A1 (n_0_115_4), .A2 (n_0_115_2), .A3 (n_0_115_6));
NAND3_X1 i_0_115_23 (.ZN (n_0_115_22), .A1 (n_0_115_1), .A2 (n_0_115_3), .A3 (n_0_115_5));
NAND3_X1 i_0_115_22 (.ZN (n_0_115_21), .A1 (n_0_115_10), .A2 (n_0_115_8), .A3 (n_0_115_12));
NAND3_X1 i_0_115_21 (.ZN (n_0_115_20), .A1 (n_0_115_7), .A2 (n_0_115_9), .A3 (n_0_115_11));
NAND2_X1 i_0_115_20 (.ZN (n_0_115_19), .A1 (n_0_115_30), .A2 (\mem[6][2] ));
INV_X1 i_0_115_19 (.ZN (n_0_115_18), .A (sps__n99));
NAND4_X1 i_0_115_18 (.ZN (n_0_115_17), .A1 (n_0_115_18), .A2 (sps__n3), .A3 (sps__n121), .A4 (sps__n112));
INV_X1 i_0_115_17 (.ZN (n_0_115_16), .A (sps__n19));
INV_X1 i_0_115_16 (.ZN (n_0_115_15), .A (sps__n81));
INV_X1 i_0_115_15 (.ZN (n_0_115_14), .A (sps__n104));
NAND3_X1 i_0_115_14 (.ZN (n_0_115_13), .A1 (n_0_115_16), .A2 (n_0_115_15), .A3 (n_0_115_14));
INV_X1 i_0_115_13 (.ZN (n_0_115_12), .A (sps__n63));
INV_X1 i_0_115_12 (.ZN (n_0_115_11), .A (sps__n75));
INV_X1 i_0_115_11 (.ZN (n_0_115_10), .A (sps__n8));
INV_X1 i_0_115_10 (.ZN (n_0_115_9), .A (sps__n14));
INV_X1 i_0_115_9 (.ZN (n_0_115_8), .A (sps__n87));
INV_X1 i_0_115_8 (.ZN (n_0_115_7), .A (sps__n34));
INV_X1 i_0_115_7 (.ZN (n_0_115_6), .A (sps__n91));
INV_X1 i_0_115_6 (.ZN (n_0_115_5), .A (sps__n67));
INV_X1 i_0_115_5 (.ZN (n_0_115_4), .A (sps__n27));
INV_X1 i_0_115_4 (.ZN (n_0_115_3), .A (sps__n44));
INV_X1 i_0_115_3 (.ZN (n_0_115_2), .A (sps__n50));
INV_X1 i_0_115_2 (.ZN (n_0_115_1), .A (sps__n57));
NAND4_X1 i_0_115_1 (.ZN (n_0_115_0), .A1 (n_0_115_26), .A2 (n_0_115_25), .A3 (n_0_115_24), .A4 (data[2]));
NAND2_X1 i_0_115_0 (.ZN (n_0_1), .A1 (n_0_115_19), .A2 (n_0_115_0));
NOR2_X1 i_0_98_34 (.ZN (n_0_98_33), .A1 (n_0_98_19), .A2 (n_0_98_0));
INV_X1 i_0_98_33 (.ZN (n_0_98_32), .A (n_0_98_0));
INV_X1 i_0_98_28 (.ZN (n_0_98_31), .A (n_0_98_19));
NAND2_X1 i_0_98_27 (.ZN (n_0_98_30), .A1 (n_0_98_29), .A2 (\mem[9][2] ));
NAND3_X1 i_0_98_23 (.ZN (n_0_98_29), .A1 (n_0_98_5), .A2 (n_0_98_32), .A3 (n_0_98_10));
NAND3_X1 i_0_98_22 (.ZN (n_0_98_28), .A1 (n_0_98_27), .A2 (n_0_98_33), .A3 (n_0_98_14));
NOR2_X1 i_0_98_21 (.ZN (n_0_98_27), .A1 (n_0_98_6), .A2 (n_0_98_26));
NAND2_X1 i_0_98_20 (.ZN (n_0_98_26), .A1 (n_0_98_10), .A2 (data[2]));
NAND2_X1 i_0_98_19 (.ZN (n_0_98_25), .A1 (n_0_98_31), .A2 (n_0_98_14));
NAND3_X1 i_0_98_18 (.ZN (n_0_0), .A1 (n_0_98_28), .A2 (n_0_98_30), .A3 (n_0_98_24));
NAND2_X1 i_0_98_17 (.ZN (n_0_98_24), .A1 (n_0_98_25), .A2 (\mem[9][2] ));
INV_X1 i_0_98_32 (.ZN (n_0_98_23), .A (sps__n34));
INV_X1 i_0_98_31 (.ZN (n_0_98_22), .A (sps__n8));
INV_X1 i_0_98_30 (.ZN (n_0_98_21), .A (sps__n14));
INV_X1 i_0_98_29 (.ZN (n_0_98_20), .A (sps__n50));
NAND4_X1 i_0_98_3 (.ZN (n_0_98_19), .A1 (n_0_98_23), .A2 (n_0_98_22), .A3 (n_0_98_21), .A4 (n_0_98_20));
INV_X1 i_0_98_26 (.ZN (n_0_98_18), .A (sps__n63));
INV_X1 i_0_98_25 (.ZN (n_0_98_17), .A (sps__n75));
INV_X1 i_0_98_24 (.ZN (n_0_98_16), .A (sps__n87));
NAND4_X1 i_0_98_6 (.ZN (n_0_98_15), .A1 (n_0_98_18), .A2 (n_0_98_17), .A3 (n_0_98_16), .A4 (sps__n1));
INV_X1 i_0_98_16 (.ZN (n_0_98_14), .A (n_0_98_15));
INV_X1 i_0_98_15 (.ZN (n_0_98_13), .A (sps__n121));
INV_X1 i_0_98_14 (.ZN (n_0_98_12), .A (sps__n112));
NAND3_X1 i_0_98_13 (.ZN (n_0_98_11), .A1 (n_0_98_13), .A2 (n_0_98_12), .A3 (sps__n97));
INV_X1 i_0_98_12 (.ZN (n_0_98_10), .A (n_0_98_11));
INV_X1 i_0_98_11 (.ZN (n_0_98_9), .A (sps__n67));
INV_X1 i_0_98_10 (.ZN (n_0_98_8), .A (sps__n19));
INV_X1 i_0_98_9 (.ZN (n_0_98_7), .A (sps__n80));
NAND4_X1 i_0_98_8 (.ZN (n_0_98_6), .A1 (n_0_98_9), .A2 (n_0_98_8), .A3 (n_0_98_7), .A4 (sps__n104));
INV_X1 i_0_98_7 (.ZN (n_0_98_5), .A (n_0_98_6));
INV_X1 i_0_98_5 (.ZN (n_0_98_4), .A (sps__n57));
INV_X1 i_0_98_4 (.ZN (n_0_98_3), .A (sps__n27));
INV_X1 i_0_98_2 (.ZN (n_0_98_2), .A (sps__n44));
INV_X1 i_0_98_1 (.ZN (n_0_98_1), .A (sps__n91));
NAND4_X1 i_0_98_0 (.ZN (n_0_98_0), .A1 (n_0_98_4), .A2 (n_0_98_3), .A3 (n_0_98_2), .A4 (n_0_98_1));
NOR2_X1 i_0_47_34 (.ZN (n_0_47_33), .A1 (n_0_47_19), .A2 (n_0_47_0));
INV_X1 i_0_47_33 (.ZN (n_0_47_32), .A (n_0_47_0));
INV_X1 i_0_47_28 (.ZN (n_0_47_31), .A (n_0_47_19));
NAND2_X1 i_0_47_27 (.ZN (n_0_47_30), .A1 (n_0_47_29), .A2 (\mem[10][2] ));
NAND3_X1 i_0_47_23 (.ZN (n_0_47_29), .A1 (n_0_47_5), .A2 (n_0_47_32), .A3 (n_0_47_10));
NAND3_X1 i_0_47_22 (.ZN (n_0_47_28), .A1 (n_0_47_27), .A2 (n_0_47_33), .A3 (n_0_47_14));
NOR2_X1 i_0_47_21 (.ZN (n_0_47_27), .A1 (n_0_47_6), .A2 (n_0_47_26));
NAND2_X1 i_0_47_20 (.ZN (n_0_47_26), .A1 (n_0_47_10), .A2 (data[2]));
NAND2_X1 i_0_47_19 (.ZN (n_0_47_25), .A1 (n_0_47_31), .A2 (n_0_47_14));
NAND3_X1 i_0_47_18 (.ZN (n_0_198), .A1 (n_0_47_28), .A2 (n_0_47_30), .A3 (n_0_47_24));
NAND2_X1 i_0_47_17 (.ZN (n_0_47_24), .A1 (n_0_47_25), .A2 (\mem[10][2] ));
INV_X1 i_0_47_32 (.ZN (n_0_47_23), .A (sps__n35));
INV_X1 i_0_47_31 (.ZN (n_0_47_22), .A (sps__n8));
INV_X1 i_0_47_30 (.ZN (n_0_47_21), .A (sps__n13));
INV_X1 i_0_47_29 (.ZN (n_0_47_20), .A (sps__n50));
NAND4_X1 i_0_47_3 (.ZN (n_0_47_19), .A1 (n_0_47_23), .A2 (n_0_47_22), .A3 (n_0_47_21), .A4 (n_0_47_20));
INV_X1 i_0_47_26 (.ZN (n_0_47_18), .A (sps__n63));
INV_X1 i_0_47_25 (.ZN (n_0_47_17), .A (sps__n75));
INV_X1 i_0_47_24 (.ZN (n_0_47_16), .A (sps__n87));
NAND4_X1 i_0_47_6 (.ZN (n_0_47_15), .A1 (n_0_47_18), .A2 (n_0_47_17), .A3 (n_0_47_16), .A4 (sps__n1));
INV_X1 i_0_47_16 (.ZN (n_0_47_14), .A (n_0_47_15));
INV_X1 i_0_47_15 (.ZN (n_0_47_13), .A (sps__n121));
INV_X1 i_0_47_14 (.ZN (n_0_47_12), .A (sps__n97));
NAND3_X1 i_0_47_13 (.ZN (n_0_47_11), .A1 (n_0_47_13), .A2 (n_0_47_12), .A3 (sps__n112));
INV_X1 i_0_47_12 (.ZN (n_0_47_10), .A (n_0_47_11));
INV_X1 i_0_47_11 (.ZN (n_0_47_9), .A (sps__n67));
INV_X1 i_0_47_10 (.ZN (n_0_47_8), .A (sps__n21));
INV_X1 i_0_47_9 (.ZN (n_0_47_7), .A (sps__n80));
NAND4_X1 i_0_47_8 (.ZN (n_0_47_6), .A1 (n_0_47_9), .A2 (n_0_47_8), .A3 (n_0_47_7), .A4 (sps__n103));
INV_X1 i_0_47_7 (.ZN (n_0_47_5), .A (n_0_47_6));
INV_X1 i_0_47_5 (.ZN (n_0_47_4), .A (sps__n57));
INV_X1 i_0_47_4 (.ZN (n_0_47_3), .A (sps__n27));
INV_X1 i_0_47_2 (.ZN (n_0_47_2), .A (sps__n44));
INV_X1 i_0_47_1 (.ZN (n_0_47_1), .A (sps__n91));
NAND4_X1 i_0_47_0 (.ZN (n_0_47_0), .A1 (n_0_47_4), .A2 (n_0_47_3), .A3 (n_0_47_2), .A4 (n_0_47_1));
NAND3_X1 i_0_30_36 (.ZN (n_0_197), .A1 (n_0_30_33), .A2 (n_0_30_34), .A3 (n_0_30_35));
NAND2_X1 i_0_30_35 (.ZN (n_0_30_35), .A1 (n_0_30_24), .A2 (\mem[1][0] ));
NAND2_X1 i_0_30_34 (.ZN (n_0_30_34), .A1 (n_0_30_23), .A2 (\mem[1][0] ));
NAND3_X1 i_0_30_33 (.ZN (n_0_30_33), .A1 (n_0_30_26), .A2 (n_0_30_32), .A3 (n_0_30_29));
NOR2_X1 i_0_30_32 (.ZN (n_0_30_32), .A1 (n_0_30_0), .A2 (n_0_30_18));
INV_X1 i_0_30_31 (.ZN (n_0_30_31), .A (n_0_30_18));
INV_X1 i_0_30_30 (.ZN (n_0_30_30), .A (n_0_30_0));
NOR2_X1 i_0_30_29 (.ZN (n_0_30_29), .A1 (n_0_30_5), .A2 (n_0_30_14));
INV_X1 i_0_30_28 (.ZN (n_0_30_28), .A (n_0_30_14));
INV_X1 i_0_30_27 (.ZN (n_0_30_27), .A (n_0_30_5));
INV_X1 i_0_30_26 (.ZN (n_0_30_26), .A (n_0_30_25));
NAND2_X1 i_0_30_25 (.ZN (n_0_30_25), .A1 (n_0_30_10), .A2 (data[0]));
NAND2_X1 i_0_30_24 (.ZN (n_0_30_24), .A1 (n_0_30_30), .A2 (n_0_30_27));
NAND3_X1 i_0_30_23 (.ZN (n_0_30_23), .A1 (n_0_30_31), .A2 (n_0_30_28), .A3 (n_0_30_10));
INV_X1 i_0_30_22 (.ZN (n_0_30_22), .A (sps__n35));
INV_X1 i_0_30_21 (.ZN (n_0_30_21), .A (sps__n8));
INV_X1 i_0_30_20 (.ZN (n_0_30_20), .A (sps__n13));
INV_X1 i_0_30_19 (.ZN (n_0_30_19), .A (sps__n49));
NAND4_X1 i_0_30_18 (.ZN (n_0_30_18), .A1 (n_0_30_22), .A2 (n_0_30_21), .A3 (n_0_30_20), .A4 (n_0_30_19));
INV_X1 i_0_30_17 (.ZN (n_0_30_17), .A (sps__n63));
INV_X1 i_0_30_12 (.ZN (n_0_30_16), .A (sps__n75));
INV_X1 i_0_30_11 (.ZN (n_0_30_15), .A (sps__n87));
NAND4_X1 i_0_30_6 (.ZN (n_0_30_14), .A1 (n_0_30_17), .A2 (n_0_30_16), .A3 (n_0_30_15), .A4 (sps__n1));
INV_X1 i_0_30_5 (.ZN (n_0_30_13), .A (sps__n121));
INV_X1 i_0_30_4 (.ZN (n_0_30_12), .A (sps__n112));
NAND3_X1 i_0_30_1 (.ZN (n_0_30_11), .A1 (n_0_30_13), .A2 (n_0_30_12), .A3 (sps__n97));
INV_X1 i_0_30_0 (.ZN (n_0_30_10), .A (n_0_30_11));
INV_X1 i_0_30_16 (.ZN (n_0_30_9), .A (sps__n67));
INV_X1 i_0_30_15 (.ZN (n_0_30_8), .A (sps__n21));
INV_X1 i_0_30_14 (.ZN (n_0_30_7), .A (sps__n80));
INV_X1 i_0_30_13 (.ZN (n_0_30_6), .A (sps__n106));
NAND4_X1 i_0_30_3 (.ZN (n_0_30_5), .A1 (n_0_30_9), .A2 (n_0_30_8), .A3 (n_0_30_7), .A4 (n_0_30_6));
INV_X1 i_0_30_10 (.ZN (n_0_30_4), .A (sps__n57));
INV_X1 i_0_30_9 (.ZN (n_0_30_3), .A (sps__n27));
INV_X1 i_0_30_8 (.ZN (n_0_30_2), .A (sps__n44));
INV_X1 i_0_30_7 (.ZN (n_0_30_1), .A (sps__n93));
NAND4_X1 i_0_30_2 (.ZN (n_0_30_0), .A1 (n_0_30_4), .A2 (n_0_30_3), .A3 (n_0_30_2), .A4 (n_0_30_1));
NAND3_X1 i_0_185_36 (.ZN (n_0_196), .A1 (n_0_185_33), .A2 (n_0_185_34), .A3 (n_0_185_35));
NAND2_X1 i_0_185_35 (.ZN (n_0_185_35), .A1 (n_0_185_24), .A2 (\mem[2][0] ));
NAND2_X1 i_0_185_34 (.ZN (n_0_185_34), .A1 (n_0_185_23), .A2 (\mem[2][0] ));
NAND3_X1 i_0_185_33 (.ZN (n_0_185_33), .A1 (n_0_185_26), .A2 (n_0_185_32), .A3 (n_0_185_29));
NOR2_X1 i_0_185_32 (.ZN (n_0_185_32), .A1 (n_0_185_0), .A2 (n_0_185_18));
INV_X1 i_0_185_31 (.ZN (n_0_185_31), .A (n_0_185_18));
INV_X1 i_0_185_30 (.ZN (n_0_185_30), .A (n_0_185_0));
NOR2_X1 i_0_185_29 (.ZN (n_0_185_29), .A1 (n_0_185_5), .A2 (n_0_185_14));
INV_X1 i_0_185_28 (.ZN (n_0_185_28), .A (n_0_185_14));
INV_X1 i_0_185_27 (.ZN (n_0_185_27), .A (n_0_185_5));
INV_X1 i_0_185_26 (.ZN (n_0_185_26), .A (n_0_185_25));
NAND2_X1 i_0_185_25 (.ZN (n_0_185_25), .A1 (n_0_185_10), .A2 (data[0]));
NAND2_X1 i_0_185_24 (.ZN (n_0_185_24), .A1 (n_0_185_30), .A2 (n_0_185_27));
NAND3_X1 i_0_185_23 (.ZN (n_0_185_23), .A1 (n_0_185_31), .A2 (n_0_185_28), .A3 (n_0_185_10));
INV_X1 i_0_185_22 (.ZN (n_0_185_22), .A (sps__n35));
INV_X1 i_0_185_21 (.ZN (n_0_185_21), .A (sps__n8));
INV_X1 i_0_185_20 (.ZN (n_0_185_20), .A (sps__n13));
INV_X1 i_0_185_19 (.ZN (n_0_185_19), .A (sps__n49));
NAND4_X1 i_0_185_18 (.ZN (n_0_185_18), .A1 (n_0_185_22), .A2 (n_0_185_21), .A3 (n_0_185_20), .A4 (n_0_185_19));
INV_X1 i_0_185_17 (.ZN (n_0_185_17), .A (sps__n61));
INV_X1 i_0_185_12 (.ZN (n_0_185_16), .A (sps__n73));
INV_X1 i_0_185_11 (.ZN (n_0_185_15), .A (sps__n85));
NAND4_X1 i_0_185_6 (.ZN (n_0_185_14), .A1 (n_0_185_17), .A2 (n_0_185_16), .A3 (n_0_185_15), .A4 (sps__n1));
INV_X1 i_0_185_5 (.ZN (n_0_185_13), .A (sps__n119));
INV_X1 i_0_185_4 (.ZN (n_0_185_12), .A (sps__n97));
NAND3_X1 i_0_185_1 (.ZN (n_0_185_11), .A1 (n_0_185_13), .A2 (n_0_185_12), .A3 (sps__n112));
INV_X1 i_0_185_0 (.ZN (n_0_185_10), .A (n_0_185_11));
INV_X1 i_0_185_16 (.ZN (n_0_185_9), .A (sps__n67));
INV_X1 i_0_185_15 (.ZN (n_0_185_8), .A (sps__n21));
INV_X1 i_0_185_14 (.ZN (n_0_185_7), .A (sps__n79));
INV_X1 i_0_185_13 (.ZN (n_0_185_6), .A (sps__n106));
NAND4_X1 i_0_185_3 (.ZN (n_0_185_5), .A1 (n_0_185_9), .A2 (n_0_185_8), .A3 (n_0_185_7), .A4 (n_0_185_6));
INV_X1 i_0_185_10 (.ZN (n_0_185_4), .A (sps__n57));
INV_X1 i_0_185_9 (.ZN (n_0_185_3), .A (sps__n27));
INV_X1 i_0_185_8 (.ZN (n_0_185_2), .A (sps__n44));
INV_X1 i_0_185_7 (.ZN (n_0_185_1), .A (sps__n93));
NAND4_X1 i_0_185_2 (.ZN (n_0_185_0), .A1 (n_0_185_4), .A2 (n_0_185_3), .A3 (n_0_185_2), .A4 (n_0_185_1));
NAND3_X1 i_0_168_36 (.ZN (n_0_195), .A1 (n_0_168_33), .A2 (n_0_168_34), .A3 (n_0_168_35));
NAND2_X1 i_0_168_35 (.ZN (n_0_168_35), .A1 (n_0_168_24), .A2 (\mem[4][0] ));
NAND2_X1 i_0_168_34 (.ZN (n_0_168_34), .A1 (n_0_168_23), .A2 (\mem[4][0] ));
NAND3_X1 i_0_168_33 (.ZN (n_0_168_33), .A1 (n_0_168_26), .A2 (n_0_168_32), .A3 (n_0_168_29));
NOR2_X1 i_0_168_32 (.ZN (n_0_168_32), .A1 (n_0_168_0), .A2 (n_0_168_18));
INV_X1 i_0_168_31 (.ZN (n_0_168_31), .A (n_0_168_18));
INV_X1 i_0_168_30 (.ZN (n_0_168_30), .A (n_0_168_0));
NOR2_X1 i_0_168_29 (.ZN (n_0_168_29), .A1 (n_0_168_5), .A2 (n_0_168_14));
INV_X1 i_0_168_28 (.ZN (n_0_168_28), .A (n_0_168_14));
INV_X1 i_0_168_27 (.ZN (n_0_168_27), .A (n_0_168_5));
INV_X1 i_0_168_26 (.ZN (n_0_168_26), .A (n_0_168_25));
NAND2_X1 i_0_168_25 (.ZN (n_0_168_25), .A1 (n_0_168_10), .A2 (data[0]));
NAND2_X1 i_0_168_24 (.ZN (n_0_168_24), .A1 (n_0_168_30), .A2 (n_0_168_27));
NAND3_X1 i_0_168_23 (.ZN (n_0_168_23), .A1 (n_0_168_31), .A2 (n_0_168_28), .A3 (n_0_168_10));
INV_X1 i_0_168_22 (.ZN (n_0_168_22), .A (sps__n35));
INV_X1 i_0_168_21 (.ZN (n_0_168_21), .A (sps__n8));
INV_X1 i_0_168_20 (.ZN (n_0_168_20), .A (sps__n13));
INV_X1 i_0_168_19 (.ZN (n_0_168_19), .A (sps__n49));
NAND4_X1 i_0_168_18 (.ZN (n_0_168_18), .A1 (n_0_168_22), .A2 (n_0_168_21), .A3 (n_0_168_20), .A4 (n_0_168_19));
INV_X1 i_0_168_17 (.ZN (n_0_168_17), .A (sps__n61));
INV_X1 i_0_168_12 (.ZN (n_0_168_16), .A (sps__n73));
INV_X1 i_0_168_11 (.ZN (n_0_168_15), .A (sps__n85));
NAND4_X1 i_0_168_6 (.ZN (n_0_168_14), .A1 (n_0_168_17), .A2 (n_0_168_16), .A3 (n_0_168_15), .A4 (sps__n1));
INV_X1 i_0_168_5 (.ZN (n_0_168_13), .A (sps__n112));
INV_X1 i_0_168_4 (.ZN (n_0_168_12), .A (sps__n97));
NAND3_X1 i_0_168_1 (.ZN (n_0_168_11), .A1 (n_0_168_13), .A2 (n_0_168_12), .A3 (sps__n119));
INV_X1 i_0_168_0 (.ZN (n_0_168_10), .A (n_0_168_11));
INV_X1 i_0_168_16 (.ZN (n_0_168_9), .A (sps__n67));
INV_X1 i_0_168_15 (.ZN (n_0_168_8), .A (sps__n21));
INV_X1 i_0_168_14 (.ZN (n_0_168_7), .A (sps__n79));
INV_X1 i_0_168_13 (.ZN (n_0_168_6), .A (sps__n106));
NAND4_X1 i_0_168_3 (.ZN (n_0_168_5), .A1 (n_0_168_9), .A2 (n_0_168_8), .A3 (n_0_168_7), .A4 (n_0_168_6));
INV_X1 i_0_168_10 (.ZN (n_0_168_4), .A (sps__n57));
INV_X1 i_0_168_9 (.ZN (n_0_168_3), .A (sps__n27));
INV_X1 i_0_168_8 (.ZN (n_0_168_2), .A (sps__n44));
INV_X1 i_0_168_7 (.ZN (n_0_168_1), .A (sps__n93));
NAND4_X1 i_0_168_2 (.ZN (n_0_168_0), .A1 (n_0_168_4), .A2 (n_0_168_3), .A3 (n_0_168_2), .A4 (n_0_168_1));
NAND3_X1 i_0_186_27 (.ZN (n_0_186_26), .A1 (n_0_186_23), .A2 (n_0_186_24), .A3 (n_0_186_25));
INV_X1 i_0_186_26 (.ZN (n_0_186_25), .A (n_0_186_17));
NOR2_X1 i_0_186_25 (.ZN (n_0_186_24), .A1 (n_0_186_18), .A2 (n_0_186_13));
INV_X1 i_0_186_24 (.ZN (n_0_186_23), .A (n_0_186_14));
OAI21_X1 i_0_186_23 (.ZN (n_0_186_22), .A (\mem[7][0] ), .B1 (n_0_186_12), .B2 (n_0_186_26));
NOR2_X1 i_0_186_22 (.ZN (n_0_186_21), .A1 (n_0_186_14), .A2 (n_0_186_13));
INV_X1 i_0_186_21 (.ZN (n_0_186_20), .A (n_0_186_12));
NOR2_X1 i_0_186_20 (.ZN (n_0_186_19), .A1 (n_0_186_17), .A2 (n_0_186_18));
NAND3_X1 i_0_186_19 (.ZN (n_0_186_18), .A1 (n_0_186_9), .A2 (n_0_186_7), .A3 (n_0_186_11));
NAND3_X1 i_0_186_18 (.ZN (n_0_186_17), .A1 (n_0_186_6), .A2 (n_0_186_8), .A3 (n_0_186_10));
NOR2_X1 i_0_186_17 (.ZN (n_0_186_16), .A1 (sps__n7), .A2 (sps__n13));
NOR2_X1 i_0_186_16 (.ZN (n_0_186_15), .A1 (sps__n85), .A2 (sps__n34));
NAND4_X1 i_0_186_15 (.ZN (n_0_186_14), .A1 (sps__n1), .A2 (sps__n119), .A3 (sps__n113), .A4 (sps__n97));
INV_X1 i_0_186_14 (.ZN (n_0_186_5), .A (sps__n21));
INV_X1 i_0_186_13 (.ZN (n_0_186_4), .A (sps__n79));
INV_X1 i_0_186_12 (.ZN (n_0_186_3), .A (sps__n106));
NAND3_X1 i_0_186_11 (.ZN (n_0_186_13), .A1 (n_0_186_5), .A2 (n_0_186_4), .A3 (n_0_186_3));
INV_X1 i_0_186_31 (.ZN (n_0_186_2), .A (sps__n61));
INV_X1 i_0_186_30 (.ZN (n_0_186_1), .A (sps__n73));
NAND2_X1 i_0_186_10 (.ZN (n_0_186_28), .A1 (n_0_186_2), .A2 (n_0_186_1));
INV_X1 i_0_186_9 (.ZN (n_0_186_27), .A (n_0_186_28));
NAND3_X1 i_0_186_8 (.ZN (n_0_186_12), .A1 (n_0_186_27), .A2 (n_0_186_16), .A3 (n_0_186_15));
INV_X1 i_0_186_7 (.ZN (n_0_186_11), .A (sps__n93));
INV_X1 i_0_186_6 (.ZN (n_0_186_10), .A (sps__n67));
INV_X1 i_0_186_5 (.ZN (n_0_186_9), .A (sps__n27));
INV_X1 i_0_186_4 (.ZN (n_0_186_8), .A (sps__n41));
INV_X1 i_0_186_3 (.ZN (n_0_186_7), .A (sps__n49));
INV_X1 i_0_186_2 (.ZN (n_0_186_6), .A (sps__n56));
NAND4_X1 i_0_186_1 (.ZN (n_0_186_0), .A1 (n_0_186_21), .A2 (n_0_186_20), .A3 (n_0_186_19), .A4 (data[0]));
NAND2_X1 i_0_186_0 (.ZN (n_0_194), .A1 (n_0_186_22), .A2 (n_0_186_0));
NAND3_X1 i_0_83_31 (.ZN (n_0_83_30), .A1 (n_0_83_27), .A2 (n_0_83_28), .A3 (n_0_83_29));
NOR2_X1 i_0_83_30 (.ZN (n_0_83_29), .A1 (n_0_83_13), .A2 (n_0_83_23));
NOR2_X1 i_0_83_29 (.ZN (n_0_83_28), .A1 (n_0_83_22), .A2 (n_0_83_21));
NOR2_X1 i_0_83_28 (.ZN (n_0_83_27), .A1 (n_0_83_17), .A2 (n_0_83_20));
NOR2_X1 i_0_83_27 (.ZN (n_0_83_26), .A1 (n_0_83_17), .A2 (n_0_83_13));
NOR2_X1 i_0_83_26 (.ZN (n_0_83_25), .A1 (n_0_83_20), .A2 (n_0_83_21));
NOR2_X1 i_0_83_25 (.ZN (n_0_83_24), .A1 (n_0_83_22), .A2 (n_0_83_23));
NAND3_X1 i_0_83_24 (.ZN (n_0_83_23), .A1 (n_0_83_4), .A2 (n_0_83_2), .A3 (n_0_83_6));
NAND3_X1 i_0_83_23 (.ZN (n_0_83_22), .A1 (n_0_83_1), .A2 (n_0_83_3), .A3 (n_0_83_5));
NAND3_X1 i_0_83_22 (.ZN (n_0_83_21), .A1 (n_0_83_10), .A2 (n_0_83_8), .A3 (n_0_83_12));
NAND3_X1 i_0_83_21 (.ZN (n_0_83_20), .A1 (n_0_83_7), .A2 (n_0_83_9), .A3 (n_0_83_11));
NAND2_X1 i_0_83_20 (.ZN (n_0_83_19), .A1 (n_0_83_30), .A2 (\mem[3][3] ));
INV_X1 i_0_83_19 (.ZN (n_0_83_18), .A (sps__n121));
NAND4_X1 i_0_83_18 (.ZN (n_0_83_17), .A1 (n_0_83_18), .A2 (sps__n1), .A3 (sps__n114), .A4 (sps__n97));
INV_X1 i_0_83_17 (.ZN (n_0_83_16), .A (sps__n21));
INV_X1 i_0_83_16 (.ZN (n_0_83_15), .A (sps__n80));
INV_X1 i_0_83_15 (.ZN (n_0_83_14), .A (sps__n103));
NAND3_X1 i_0_83_14 (.ZN (n_0_83_13), .A1 (n_0_83_16), .A2 (n_0_83_15), .A3 (n_0_83_14));
INV_X1 i_0_83_13 (.ZN (n_0_83_12), .A (sps__n61));
INV_X1 i_0_83_12 (.ZN (n_0_83_11), .A (sps__n74));
INV_X1 i_0_83_11 (.ZN (n_0_83_10), .A (sps__n7));
INV_X1 i_0_83_10 (.ZN (n_0_83_9), .A (address[12]));
INV_X1 i_0_83_9 (.ZN (n_0_83_8), .A (sps__n87));
INV_X1 i_0_83_8 (.ZN (n_0_83_7), .A (sps__n36));
INV_X1 i_0_83_7 (.ZN (n_0_83_6), .A (sps__n91));
INV_X1 i_0_83_6 (.ZN (n_0_83_5), .A (sps__n69));
INV_X1 i_0_83_5 (.ZN (n_0_83_4), .A (sps__n27));
INV_X1 i_0_83_4 (.ZN (n_0_83_3), .A (sps__n41));
INV_X1 i_0_83_3 (.ZN (n_0_83_2), .A (sps__n49));
INV_X1 i_0_83_2 (.ZN (n_0_83_1), .A (sps__n56));
NAND4_X1 i_0_83_1 (.ZN (n_0_83_0), .A1 (n_0_83_26), .A2 (n_0_83_25), .A3 (n_0_83_24), .A4 (data[3]));
NAND2_X1 i_0_83_0 (.ZN (n_0_193), .A1 (n_0_83_19), .A2 (n_0_83_0));
NAND3_X1 i_0_148_31 (.ZN (n_0_148_30), .A1 (n_0_148_27), .A2 (n_0_148_28), .A3 (n_0_148_29));
NOR2_X1 i_0_148_30 (.ZN (n_0_148_29), .A1 (n_0_148_13), .A2 (n_0_148_23));
NOR2_X1 i_0_148_29 (.ZN (n_0_148_28), .A1 (n_0_148_22), .A2 (n_0_148_21));
NOR2_X1 i_0_148_28 (.ZN (n_0_148_27), .A1 (n_0_148_17), .A2 (n_0_148_20));
NOR2_X1 i_0_148_27 (.ZN (n_0_148_26), .A1 (n_0_148_17), .A2 (n_0_148_13));
NOR2_X1 i_0_148_26 (.ZN (n_0_148_25), .A1 (n_0_148_20), .A2 (n_0_148_21));
NOR2_X1 i_0_148_25 (.ZN (n_0_148_24), .A1 (n_0_148_22), .A2 (n_0_148_23));
NAND3_X1 i_0_148_24 (.ZN (n_0_148_23), .A1 (n_0_148_4), .A2 (n_0_148_2), .A3 (n_0_148_6));
NAND3_X1 i_0_148_23 (.ZN (n_0_148_22), .A1 (n_0_148_1), .A2 (n_0_148_3), .A3 (n_0_148_5));
NAND3_X1 i_0_148_22 (.ZN (n_0_148_21), .A1 (n_0_148_10), .A2 (n_0_148_8), .A3 (n_0_148_12));
NAND3_X1 i_0_148_21 (.ZN (n_0_148_20), .A1 (n_0_148_7), .A2 (n_0_148_9), .A3 (n_0_148_11));
NAND2_X1 i_0_148_20 (.ZN (n_0_148_19), .A1 (n_0_148_30), .A2 (\mem[5][3] ));
INV_X1 i_0_148_19 (.ZN (n_0_148_18), .A (sps__n112));
NAND4_X1 i_0_148_18 (.ZN (n_0_148_17), .A1 (n_0_148_18), .A2 (sps__n3), .A3 (sps__n121), .A4 (sps__n99));
INV_X1 i_0_148_17 (.ZN (n_0_148_16), .A (sps__n21));
INV_X1 i_0_148_16 (.ZN (n_0_148_15), .A (sps__n80));
INV_X1 i_0_148_15 (.ZN (n_0_148_14), .A (sps__n103));
NAND3_X1 i_0_148_14 (.ZN (n_0_148_13), .A1 (n_0_148_16), .A2 (n_0_148_15), .A3 (n_0_148_14));
INV_X1 i_0_148_13 (.ZN (n_0_148_12), .A (sps__n62));
INV_X1 i_0_148_12 (.ZN (n_0_148_11), .A (sps__n74));
INV_X1 i_0_148_11 (.ZN (n_0_148_10), .A (sps__n8));
INV_X1 i_0_148_10 (.ZN (n_0_148_9), .A (sps__n14));
INV_X1 i_0_148_9 (.ZN (n_0_148_8), .A (sps__n85));
INV_X1 i_0_148_8 (.ZN (n_0_148_7), .A (sps__n34));
INV_X1 i_0_148_7 (.ZN (n_0_148_6), .A (sps__n91));
INV_X1 i_0_148_6 (.ZN (n_0_148_5), .A (sps__n68));
INV_X1 i_0_148_5 (.ZN (n_0_148_4), .A (sps__n26));
INV_X1 i_0_148_4 (.ZN (n_0_148_3), .A (sps__n44));
INV_X1 i_0_148_3 (.ZN (n_0_148_2), .A (sps__n49));
INV_X1 i_0_148_2 (.ZN (n_0_148_1), .A (sps__n55));
NAND4_X1 i_0_148_1 (.ZN (n_0_148_0), .A1 (n_0_148_26), .A2 (n_0_148_25), .A3 (n_0_148_24), .A4 (data[3]));
NAND2_X1 i_0_148_0 (.ZN (n_0_192), .A1 (n_0_148_19), .A2 (n_0_148_0));
NAND3_X1 i_0_114_31 (.ZN (n_0_114_30), .A1 (n_0_114_27), .A2 (n_0_114_28), .A3 (n_0_114_29));
NOR2_X1 i_0_114_30 (.ZN (n_0_114_29), .A1 (n_0_114_13), .A2 (n_0_114_23));
NOR2_X1 i_0_114_29 (.ZN (n_0_114_28), .A1 (n_0_114_22), .A2 (n_0_114_21));
NOR2_X1 i_0_114_28 (.ZN (n_0_114_27), .A1 (n_0_114_17), .A2 (n_0_114_20));
NOR2_X1 i_0_114_27 (.ZN (n_0_114_26), .A1 (n_0_114_17), .A2 (n_0_114_13));
NOR2_X1 i_0_114_26 (.ZN (n_0_114_25), .A1 (n_0_114_20), .A2 (n_0_114_21));
NOR2_X1 i_0_114_25 (.ZN (n_0_114_24), .A1 (n_0_114_22), .A2 (n_0_114_23));
NAND3_X1 i_0_114_24 (.ZN (n_0_114_23), .A1 (n_0_114_4), .A2 (n_0_114_2), .A3 (n_0_114_6));
NAND3_X1 i_0_114_23 (.ZN (n_0_114_22), .A1 (n_0_114_1), .A2 (n_0_114_3), .A3 (n_0_114_5));
NAND3_X1 i_0_114_22 (.ZN (n_0_114_21), .A1 (n_0_114_10), .A2 (n_0_114_8), .A3 (n_0_114_12));
NAND3_X1 i_0_114_21 (.ZN (n_0_114_20), .A1 (n_0_114_7), .A2 (n_0_114_9), .A3 (n_0_114_11));
NAND2_X1 i_0_114_20 (.ZN (n_0_114_19), .A1 (n_0_114_30), .A2 (\mem[6][3] ));
INV_X1 i_0_114_19 (.ZN (n_0_114_18), .A (sps__n99));
NAND4_X1 i_0_114_18 (.ZN (n_0_114_17), .A1 (n_0_114_18), .A2 (sps__n3), .A3 (sps__n122), .A4 (sps__n112));
INV_X1 i_0_114_17 (.ZN (n_0_114_16), .A (sps__n19));
INV_X1 i_0_114_16 (.ZN (n_0_114_15), .A (sps__n81));
INV_X1 i_0_114_15 (.ZN (n_0_114_14), .A (sps__n105));
NAND3_X1 i_0_114_14 (.ZN (n_0_114_13), .A1 (n_0_114_16), .A2 (n_0_114_15), .A3 (n_0_114_14));
INV_X1 i_0_114_13 (.ZN (n_0_114_12), .A (sps__n62));
INV_X1 i_0_114_12 (.ZN (n_0_114_11), .A (sps__n75));
INV_X1 i_0_114_11 (.ZN (n_0_114_10), .A (sps__n9));
INV_X1 i_0_114_10 (.ZN (n_0_114_9), .A (sps__n15));
INV_X1 i_0_114_9 (.ZN (n_0_114_8), .A (sps__n86));
INV_X1 i_0_114_8 (.ZN (n_0_114_7), .A (sps__n34));
INV_X1 i_0_114_7 (.ZN (n_0_114_6), .A (sps__n92));
INV_X1 i_0_114_6 (.ZN (n_0_114_5), .A (sps__n67));
INV_X1 i_0_114_5 (.ZN (n_0_114_4), .A (sps__n28));
INV_X1 i_0_114_4 (.ZN (n_0_114_3), .A (sps__n43));
INV_X1 i_0_114_3 (.ZN (n_0_114_2), .A (sps__n51));
INV_X1 i_0_114_2 (.ZN (n_0_114_1), .A (sps__n55));
NAND4_X1 i_0_114_1 (.ZN (n_0_114_0), .A1 (n_0_114_26), .A2 (n_0_114_25), .A3 (n_0_114_24), .A4 (data[3]));
NAND2_X1 i_0_114_0 (.ZN (n_0_191), .A1 (n_0_114_19), .A2 (n_0_114_0));
NOR2_X1 i_0_97_34 (.ZN (n_0_97_33), .A1 (n_0_97_19), .A2 (n_0_97_0));
INV_X1 i_0_97_33 (.ZN (n_0_97_32), .A (n_0_97_0));
INV_X1 i_0_97_28 (.ZN (n_0_97_31), .A (n_0_97_19));
NAND2_X1 i_0_97_27 (.ZN (n_0_97_30), .A1 (n_0_97_29), .A2 (\mem[9][3] ));
NAND3_X1 i_0_97_23 (.ZN (n_0_97_29), .A1 (n_0_97_5), .A2 (n_0_97_32), .A3 (n_0_97_10));
NAND3_X1 i_0_97_22 (.ZN (n_0_97_28), .A1 (n_0_97_27), .A2 (n_0_97_33), .A3 (n_0_97_14));
NOR2_X1 i_0_97_21 (.ZN (n_0_97_27), .A1 (n_0_97_6), .A2 (n_0_97_26));
NAND2_X1 i_0_97_20 (.ZN (n_0_97_26), .A1 (n_0_97_10), .A2 (data[3]));
NAND2_X1 i_0_97_19 (.ZN (n_0_97_25), .A1 (n_0_97_31), .A2 (n_0_97_14));
NAND3_X1 i_0_97_18 (.ZN (n_0_190), .A1 (n_0_97_28), .A2 (n_0_97_30), .A3 (n_0_97_24));
NAND2_X1 i_0_97_17 (.ZN (n_0_97_24), .A1 (n_0_97_25), .A2 (\mem[9][3] ));
INV_X1 i_0_97_32 (.ZN (n_0_97_23), .A (sps__n34));
INV_X1 i_0_97_31 (.ZN (n_0_97_22), .A (sps__n8));
INV_X1 i_0_97_30 (.ZN (n_0_97_21), .A (sps__n14));
INV_X1 i_0_97_29 (.ZN (n_0_97_20), .A (sps__n50));
NAND4_X1 i_0_97_3 (.ZN (n_0_97_19), .A1 (n_0_97_23), .A2 (n_0_97_22), .A3 (n_0_97_21), .A4 (n_0_97_20));
INV_X1 i_0_97_26 (.ZN (n_0_97_18), .A (sps__n63));
INV_X1 i_0_97_25 (.ZN (n_0_97_17), .A (sps__n74));
INV_X1 i_0_97_24 (.ZN (n_0_97_16), .A (sps__n87));
NAND4_X1 i_0_97_6 (.ZN (n_0_97_15), .A1 (n_0_97_18), .A2 (n_0_97_17), .A3 (n_0_97_16), .A4 (sps__n3));
INV_X1 i_0_97_16 (.ZN (n_0_97_14), .A (n_0_97_15));
INV_X1 i_0_97_15 (.ZN (n_0_97_13), .A (sps__n122));
INV_X1 i_0_97_14 (.ZN (n_0_97_12), .A (sps__n112));
NAND3_X1 i_0_97_13 (.ZN (n_0_97_11), .A1 (n_0_97_13), .A2 (n_0_97_12), .A3 (sps__n99));
INV_X1 i_0_97_12 (.ZN (n_0_97_10), .A (n_0_97_11));
INV_X1 i_0_97_11 (.ZN (n_0_97_9), .A (sps__n68));
INV_X1 i_0_97_10 (.ZN (n_0_97_8), .A (sps__n19));
INV_X1 i_0_97_9 (.ZN (n_0_97_7), .A (sps__n81));
NAND4_X1 i_0_97_8 (.ZN (n_0_97_6), .A1 (n_0_97_9), .A2 (n_0_97_8), .A3 (n_0_97_7), .A4 (sps__n104));
INV_X1 i_0_97_7 (.ZN (n_0_97_5), .A (n_0_97_6));
INV_X1 i_0_97_5 (.ZN (n_0_97_4), .A (sps__n57));
INV_X1 i_0_97_4 (.ZN (n_0_97_3), .A (sps__n26));
INV_X1 i_0_97_2 (.ZN (n_0_97_2), .A (sps__n44));
INV_X1 i_0_97_1 (.ZN (n_0_97_1), .A (sps__n91));
NAND4_X1 i_0_97_0 (.ZN (n_0_97_0), .A1 (n_0_97_4), .A2 (n_0_97_3), .A3 (n_0_97_2), .A4 (n_0_97_1));
NOR2_X1 i_0_46_34 (.ZN (n_0_46_33), .A1 (n_0_46_19), .A2 (n_0_46_0));
INV_X1 i_0_46_33 (.ZN (n_0_46_32), .A (n_0_46_0));
INV_X1 i_0_46_28 (.ZN (n_0_46_31), .A (n_0_46_19));
NAND2_X1 i_0_46_27 (.ZN (n_0_46_30), .A1 (n_0_46_29), .A2 (\mem[10][3] ));
NAND3_X1 i_0_46_23 (.ZN (n_0_46_29), .A1 (n_0_46_5), .A2 (n_0_46_32), .A3 (n_0_46_10));
NAND3_X1 i_0_46_22 (.ZN (n_0_46_28), .A1 (n_0_46_27), .A2 (n_0_46_33), .A3 (n_0_46_14));
NOR2_X1 i_0_46_21 (.ZN (n_0_46_27), .A1 (n_0_46_6), .A2 (n_0_46_26));
NAND2_X1 i_0_46_20 (.ZN (n_0_46_26), .A1 (n_0_46_10), .A2 (data[3]));
NAND2_X1 i_0_46_19 (.ZN (n_0_46_25), .A1 (n_0_46_31), .A2 (n_0_46_14));
NAND3_X1 i_0_46_18 (.ZN (n_0_189), .A1 (n_0_46_28), .A2 (n_0_46_30), .A3 (n_0_46_24));
NAND2_X1 i_0_46_17 (.ZN (n_0_46_24), .A1 (n_0_46_25), .A2 (\mem[10][3] ));
INV_X1 i_0_46_32 (.ZN (n_0_46_23), .A (sps__n34));
INV_X1 i_0_46_31 (.ZN (n_0_46_22), .A (sps__n8));
INV_X1 i_0_46_30 (.ZN (n_0_46_21), .A (sps__n14));
INV_X1 i_0_46_29 (.ZN (n_0_46_20), .A (sps__n50));
NAND4_X1 i_0_46_3 (.ZN (n_0_46_19), .A1 (n_0_46_23), .A2 (n_0_46_22), .A3 (n_0_46_21), .A4 (n_0_46_20));
INV_X1 i_0_46_26 (.ZN (n_0_46_18), .A (sps__n63));
INV_X1 i_0_46_25 (.ZN (n_0_46_17), .A (sps__n74));
INV_X1 i_0_46_24 (.ZN (n_0_46_16), .A (sps__n86));
NAND4_X1 i_0_46_6 (.ZN (n_0_46_15), .A1 (n_0_46_18), .A2 (n_0_46_17), .A3 (n_0_46_16), .A4 (sps__n3));
INV_X1 i_0_46_16 (.ZN (n_0_46_14), .A (n_0_46_15));
INV_X1 i_0_46_15 (.ZN (n_0_46_13), .A (sps__n121));
INV_X1 i_0_46_14 (.ZN (n_0_46_12), .A (sps__n99));
NAND3_X1 i_0_46_13 (.ZN (n_0_46_11), .A1 (n_0_46_13), .A2 (n_0_46_12), .A3 (sps__n112));
INV_X1 i_0_46_12 (.ZN (n_0_46_10), .A (n_0_46_11));
INV_X1 i_0_46_11 (.ZN (n_0_46_9), .A (sps__n68));
INV_X1 i_0_46_10 (.ZN (n_0_46_8), .A (sps__n19));
INV_X1 i_0_46_9 (.ZN (n_0_46_7), .A (sps__n81));
NAND4_X1 i_0_46_8 (.ZN (n_0_46_6), .A1 (n_0_46_9), .A2 (n_0_46_8), .A3 (n_0_46_7), .A4 (sps__n104));
INV_X1 i_0_46_7 (.ZN (n_0_46_5), .A (n_0_46_6));
INV_X1 i_0_46_5 (.ZN (n_0_46_4), .A (sps__n55));
INV_X1 i_0_46_4 (.ZN (n_0_46_3), .A (sps__n28));
INV_X1 i_0_46_2 (.ZN (n_0_46_2), .A (sps__n44));
INV_X1 i_0_46_1 (.ZN (n_0_46_1), .A (sps__n92));
NAND4_X1 i_0_46_0 (.ZN (n_0_46_0), .A1 (n_0_46_4), .A2 (n_0_46_3), .A3 (n_0_46_2), .A4 (n_0_46_1));
NAND3_X1 i_0_29_27 (.ZN (n_0_29_26), .A1 (n_0_29_23), .A2 (n_0_29_24), .A3 (n_0_29_25));
NOR2_X1 i_0_29_26 (.ZN (n_0_29_25), .A1 (n_0_29_17), .A2 (n_0_29_13));
NOR2_X1 i_0_29_25 (.ZN (n_0_29_24), .A1 (n_0_29_19), .A2 (n_0_29_20));
NOR2_X1 i_0_29_24 (.ZN (n_0_29_23), .A1 (n_0_29_21), .A2 (n_0_29_22));
NAND3_X1 i_0_29_23 (.ZN (n_0_29_22), .A1 (n_0_29_4), .A2 (n_0_29_2), .A3 (n_0_29_6));
NAND3_X1 i_0_29_22 (.ZN (n_0_29_21), .A1 (n_0_29_1), .A2 (n_0_29_3), .A3 (n_0_29_5));
NAND3_X1 i_0_29_21 (.ZN (n_0_29_20), .A1 (n_0_29_10), .A2 (n_0_29_8), .A3 (n_0_29_12));
NAND3_X1 i_0_29_20 (.ZN (n_0_29_19), .A1 (n_0_29_7), .A2 (n_0_29_9), .A3 (n_0_29_11));
NAND2_X1 i_0_29_19 (.ZN (n_0_29_18), .A1 (n_0_29_26), .A2 (\mem[7][1] ));
NAND4_X1 i_0_29_18 (.ZN (n_0_29_17), .A1 (sps__n1), .A2 (sps__n119), .A3 (sps__n113), .A4 (address[0]));
INV_X1 i_0_29_17 (.ZN (n_0_29_16), .A (sps__n21));
INV_X1 i_0_29_16 (.ZN (n_0_29_15), .A (sps__n79));
INV_X1 i_0_29_15 (.ZN (n_0_29_14), .A (sps__n106));
NAND3_X1 i_0_29_14 (.ZN (n_0_29_13), .A1 (n_0_29_16), .A2 (n_0_29_15), .A3 (n_0_29_14));
INV_X1 i_0_29_13 (.ZN (n_0_29_12), .A (sps__n61));
INV_X1 i_0_29_12 (.ZN (n_0_29_11), .A (sps__n73));
INV_X1 i_0_29_11 (.ZN (n_0_29_10), .A (sps__n7));
INV_X1 i_0_29_10 (.ZN (n_0_29_9), .A (sps__n13));
INV_X1 i_0_29_9 (.ZN (n_0_29_8), .A (sps__n85));
INV_X1 i_0_29_8 (.ZN (n_0_29_7), .A (sps__n34));
INV_X1 i_0_29_7 (.ZN (n_0_29_6), .A (sps__n93));
INV_X1 i_0_29_6 (.ZN (n_0_29_5), .A (sps__n69));
INV_X1 i_0_29_5 (.ZN (n_0_29_4), .A (sps__n27));
INV_X1 i_0_29_4 (.ZN (n_0_29_3), .A (sps__n41));
INV_X1 i_0_29_3 (.ZN (n_0_29_2), .A (sps__n49));
INV_X1 i_0_29_2 (.ZN (n_0_29_1), .A (sps__n56));
NAND4_X1 i_0_29_1 (.ZN (n_0_29_0), .A1 (n_0_29_25), .A2 (n_0_29_24), .A3 (n_0_29_23), .A4 (data[1]));
NAND2_X1 i_0_29_0 (.ZN (n_0_188), .A1 (n_0_29_18), .A2 (n_0_29_0));
NAND3_X1 i_0_82_35 (.ZN (n_0_186), .A1 (n_0_82_32), .A2 (n_0_82_33), .A3 (n_0_82_34));
NAND2_X1 i_0_82_34 (.ZN (n_0_82_34), .A1 (n_0_82_23), .A2 (\mem[8][1] ));
NAND3_X1 i_0_82_29 (.ZN (n_0_82_33), .A1 (n_0_82_26), .A2 (n_0_82_31), .A3 (n_0_82_28));
NAND2_X1 i_0_82_28 (.ZN (n_0_82_32), .A1 (n_0_82_27), .A2 (\mem[8][1] ));
NOR2_X1 i_0_82_24 (.ZN (n_0_82_31), .A1 (n_0_82_18), .A2 (n_0_82_0));
INV_X1 i_0_82_23 (.ZN (n_0_82_30), .A (n_0_82_0));
INV_X1 i_0_82_22 (.ZN (n_0_82_29), .A (n_0_82_18));
INV_X1 i_0_82_21 (.ZN (n_0_82_28), .A (n_0_82_5));
NAND3_X1 i_0_82_20 (.ZN (n_0_82_27), .A1 (n_0_82_28), .A2 (n_0_82_30), .A3 (n_0_82_9));
NOR2_X1 i_0_82_19 (.ZN (n_0_82_26), .A1 (n_0_82_14), .A2 (n_0_82_24));
INV_X1 i_0_82_18 (.ZN (n_0_82_25), .A (n_0_82_14));
NAND2_X1 i_0_82_17 (.ZN (n_0_82_24), .A1 (n_0_82_9), .A2 (data[1]));
NAND2_X1 i_0_82_16 (.ZN (n_0_82_23), .A1 (n_0_82_29), .A2 (n_0_82_25));
INV_X1 i_0_82_33 (.ZN (n_0_82_22), .A (sps__n34));
INV_X1 i_0_82_32 (.ZN (n_0_82_21), .A (sps__n7));
INV_X1 i_0_82_31 (.ZN (n_0_82_20), .A (sps__n13));
INV_X1 i_0_82_30 (.ZN (n_0_82_19), .A (sps__n49));
NAND4_X1 i_0_82_3 (.ZN (n_0_82_18), .A1 (n_0_82_22), .A2 (n_0_82_21), .A3 (n_0_82_20), .A4 (n_0_82_19));
INV_X1 i_0_82_27 (.ZN (n_0_82_17), .A (sps__n61));
INV_X1 i_0_82_26 (.ZN (n_0_82_16), .A (sps__n73));
INV_X1 i_0_82_25 (.ZN (n_0_82_15), .A (sps__n85));
NAND4_X1 i_0_82_8 (.ZN (n_0_82_14), .A1 (n_0_82_17), .A2 (n_0_82_16), .A3 (n_0_82_15), .A4 (sps__n1));
INV_X1 i_0_82_15 (.ZN (n_0_82_13), .A (sps__n119));
INV_X1 i_0_82_14 (.ZN (n_0_82_12), .A (sps__n113));
INV_X1 i_0_82_13 (.ZN (n_0_82_11), .A (address[0]));
NAND3_X1 i_0_82_12 (.ZN (n_0_82_10), .A1 (n_0_82_13), .A2 (n_0_82_12), .A3 (n_0_82_11));
INV_X1 i_0_82_11 (.ZN (n_0_82_9), .A (n_0_82_10));
INV_X1 i_0_82_10 (.ZN (n_0_82_8), .A (sps__n69));
INV_X1 i_0_82_9 (.ZN (n_0_82_7), .A (sps__n21));
INV_X1 i_0_82_7 (.ZN (n_0_82_6), .A (sps__n79));
NAND4_X1 i_0_82_6 (.ZN (n_0_82_5), .A1 (n_0_82_8), .A2 (n_0_82_7), .A3 (n_0_82_6), .A4 (sps__n106));
INV_X1 i_0_82_5 (.ZN (n_0_82_4), .A (sps__n56));
INV_X1 i_0_82_4 (.ZN (n_0_82_3), .A (sps__n27));
INV_X1 i_0_82_2 (.ZN (n_0_82_2), .A (sps__n41));
INV_X1 i_0_82_1 (.ZN (n_0_82_1), .A (sps__n93));
NAND4_X1 i_0_82_0 (.ZN (n_0_82_0), .A1 (n_0_82_4), .A2 (n_0_82_3), .A3 (n_0_82_2), .A4 (n_0_82_1));
NAND3_X1 i_0_65_37 (.ZN (n_0_184), .A1 (n_0_65_34), .A2 (n_0_65_35), .A3 (n_0_65_36));
NAND2_X1 i_0_65_36 (.ZN (n_0_65_36), .A1 (n_0_65_25), .A2 (\mem[0][1] ));
NAND3_X1 i_0_65_35 (.ZN (n_0_65_35), .A1 (n_0_65_27), .A2 (n_0_65_33), .A3 (n_0_65_30));
NAND2_X1 i_0_65_34 (.ZN (n_0_65_34), .A1 (n_0_65_24), .A2 (\mem[0][1] ));
NOR2_X1 i_0_65_33 (.ZN (n_0_65_33), .A1 (n_0_65_0), .A2 (n_0_65_19));
INV_X1 i_0_65_32 (.ZN (n_0_65_32), .A (n_0_65_19));
INV_X1 i_0_65_31 (.ZN (n_0_65_31), .A (n_0_65_0));
NOR2_X1 i_0_65_30 (.ZN (n_0_65_30), .A1 (n_0_65_5), .A2 (n_0_65_15));
INV_X1 i_0_65_29 (.ZN (n_0_65_29), .A (n_0_65_15));
INV_X1 i_0_65_28 (.ZN (n_0_65_28), .A (n_0_65_5));
INV_X1 i_0_65_27 (.ZN (n_0_65_27), .A (n_0_65_26));
NAND2_X1 i_0_65_26 (.ZN (n_0_65_26), .A1 (n_0_65_10), .A2 (data[1]));
NAND2_X1 i_0_65_25 (.ZN (n_0_65_25), .A1 (n_0_65_31), .A2 (n_0_65_28));
NAND3_X1 i_0_65_24 (.ZN (n_0_65_24), .A1 (n_0_65_32), .A2 (n_0_65_29), .A3 (n_0_65_10));
INV_X1 i_0_65_23 (.ZN (n_0_65_23), .A (sps__n34));
INV_X1 i_0_65_22 (.ZN (n_0_65_22), .A (sps__n7));
INV_X1 i_0_65_21 (.ZN (n_0_65_21), .A (sps__n13));
INV_X1 i_0_65_20 (.ZN (n_0_65_20), .A (sps__n49));
NAND4_X1 i_0_65_19 (.ZN (n_0_65_19), .A1 (n_0_65_23), .A2 (n_0_65_22), .A3 (n_0_65_21), .A4 (n_0_65_20));
INV_X1 i_0_65_18 (.ZN (n_0_65_18), .A (sps__n61));
INV_X1 i_0_65_17 (.ZN (n_0_65_17), .A (sps__n73));
INV_X1 i_0_65_12 (.ZN (n_0_65_16), .A (sps__n85));
NAND4_X1 i_0_65_11 (.ZN (n_0_65_15), .A1 (n_0_65_18), .A2 (n_0_65_17), .A3 (n_0_65_16), .A4 (sps__n1));
INV_X1 i_0_65_6 (.ZN (n_0_65_14), .A (sps__n119));
INV_X1 i_0_65_5 (.ZN (n_0_65_13), .A (sps__n113));
INV_X1 i_0_65_4 (.ZN (n_0_65_12), .A (address[0]));
NAND3_X1 i_0_65_1 (.ZN (n_0_65_11), .A1 (n_0_65_14), .A2 (n_0_65_13), .A3 (n_0_65_12));
INV_X1 i_0_65_0 (.ZN (n_0_65_10), .A (n_0_65_11));
INV_X1 i_0_65_16 (.ZN (n_0_65_9), .A (sps__n67));
INV_X1 i_0_65_15 (.ZN (n_0_65_8), .A (sps__n21));
INV_X1 i_0_65_14 (.ZN (n_0_65_7), .A (sps__n79));
INV_X1 i_0_65_13 (.ZN (n_0_65_6), .A (sps__n106));
NAND4_X1 i_0_65_3 (.ZN (n_0_65_5), .A1 (n_0_65_9), .A2 (n_0_65_8), .A3 (n_0_65_7), .A4 (n_0_65_6));
INV_X1 i_0_65_10 (.ZN (n_0_65_4), .A (sps__n56));
INV_X1 i_0_65_9 (.ZN (n_0_65_3), .A (sps__n27));
INV_X1 i_0_65_8 (.ZN (n_0_65_2), .A (sps__n41));
INV_X1 i_0_65_7 (.ZN (n_0_65_1), .A (sps__n93));
NAND4_X1 i_0_65_2 (.ZN (n_0_65_0), .A1 (n_0_65_4), .A2 (n_0_65_3), .A3 (n_0_65_2), .A4 (n_0_65_1));
NAND3_X1 i_0_188_36 (.ZN (n_0_183), .A1 (n_0_188_33), .A2 (n_0_188_34), .A3 (n_0_188_35));
NAND2_X1 i_0_188_35 (.ZN (n_0_188_35), .A1 (n_0_188_24), .A2 (\mem[1][1] ));
NAND2_X1 i_0_188_34 (.ZN (n_0_188_34), .A1 (n_0_188_23), .A2 (\mem[1][1] ));
NAND3_X1 i_0_188_33 (.ZN (n_0_188_33), .A1 (n_0_188_26), .A2 (n_0_188_32), .A3 (n_0_188_29));
NOR2_X1 i_0_188_32 (.ZN (n_0_188_32), .A1 (n_0_188_0), .A2 (n_0_188_18));
INV_X1 i_0_188_31 (.ZN (n_0_188_31), .A (n_0_188_18));
INV_X1 i_0_188_30 (.ZN (n_0_188_30), .A (n_0_188_0));
NOR2_X1 i_0_188_29 (.ZN (n_0_188_29), .A1 (n_0_188_5), .A2 (n_0_188_14));
INV_X1 i_0_188_28 (.ZN (n_0_188_28), .A (n_0_188_14));
INV_X1 i_0_188_27 (.ZN (n_0_188_27), .A (n_0_188_5));
INV_X1 i_0_188_26 (.ZN (n_0_188_26), .A (n_0_188_25));
NAND2_X1 i_0_188_25 (.ZN (n_0_188_25), .A1 (n_0_188_10), .A2 (data[1]));
NAND2_X1 i_0_188_24 (.ZN (n_0_188_24), .A1 (n_0_188_30), .A2 (n_0_188_27));
NAND3_X1 i_0_188_23 (.ZN (n_0_188_23), .A1 (n_0_188_31), .A2 (n_0_188_28), .A3 (n_0_188_10));
INV_X1 i_0_188_22 (.ZN (n_0_188_22), .A (sps__n36));
INV_X1 i_0_188_21 (.ZN (n_0_188_21), .A (sps__n7));
INV_X1 i_0_188_20 (.ZN (n_0_188_20), .A (sps__n13));
INV_X1 i_0_188_19 (.ZN (n_0_188_19), .A (sps__n49));
NAND4_X1 i_0_188_18 (.ZN (n_0_188_18), .A1 (n_0_188_22), .A2 (n_0_188_21), .A3 (n_0_188_20), .A4 (n_0_188_19));
INV_X1 i_0_188_17 (.ZN (n_0_188_17), .A (sps__n61));
INV_X1 i_0_188_12 (.ZN (n_0_188_16), .A (sps__n73));
INV_X1 i_0_188_11 (.ZN (n_0_188_15), .A (sps__n85));
NAND4_X1 i_0_188_6 (.ZN (n_0_188_14), .A1 (n_0_188_17), .A2 (n_0_188_16), .A3 (n_0_188_15), .A4 (sps__n1));
INV_X1 i_0_188_5 (.ZN (n_0_188_13), .A (sps__n119));
INV_X1 i_0_188_4 (.ZN (n_0_188_12), .A (sps__n113));
NAND3_X1 i_0_188_1 (.ZN (n_0_188_11), .A1 (n_0_188_13), .A2 (n_0_188_12), .A3 (sps__n97));
INV_X1 i_0_188_0 (.ZN (n_0_188_10), .A (n_0_188_11));
INV_X1 i_0_188_16 (.ZN (n_0_188_9), .A (sps__n69));
INV_X1 i_0_188_15 (.ZN (n_0_188_8), .A (sps__n21));
INV_X1 i_0_188_14 (.ZN (n_0_188_7), .A (sps__n79));
INV_X1 i_0_188_13 (.ZN (n_0_188_6), .A (sps__n103));
NAND4_X1 i_0_188_3 (.ZN (n_0_188_5), .A1 (n_0_188_9), .A2 (n_0_188_8), .A3 (n_0_188_7), .A4 (n_0_188_6));
INV_X1 i_0_188_10 (.ZN (n_0_188_4), .A (sps__n56));
INV_X1 i_0_188_9 (.ZN (n_0_188_3), .A (sps__n27));
INV_X1 i_0_188_8 (.ZN (n_0_188_2), .A (sps__n41));
INV_X1 i_0_188_7 (.ZN (n_0_188_1), .A (sps__n91));
NAND4_X1 i_0_188_2 (.ZN (n_0_188_0), .A1 (n_0_188_4), .A2 (n_0_188_3), .A3 (n_0_188_2), .A4 (n_0_188_1));
NAND3_X1 i_0_184_36 (.ZN (n_0_182), .A1 (n_0_184_33), .A2 (n_0_184_34), .A3 (n_0_184_35));
NAND2_X1 i_0_184_35 (.ZN (n_0_184_35), .A1 (n_0_184_24), .A2 (\mem[2][1] ));
NAND2_X1 i_0_184_34 (.ZN (n_0_184_34), .A1 (n_0_184_23), .A2 (\mem[2][1] ));
NAND3_X1 i_0_184_33 (.ZN (n_0_184_33), .A1 (n_0_184_26), .A2 (n_0_184_32), .A3 (n_0_184_29));
NOR2_X1 i_0_184_32 (.ZN (n_0_184_32), .A1 (n_0_184_0), .A2 (n_0_184_18));
INV_X1 i_0_184_31 (.ZN (n_0_184_31), .A (n_0_184_18));
INV_X1 i_0_184_30 (.ZN (n_0_184_30), .A (n_0_184_0));
NOR2_X1 i_0_184_29 (.ZN (n_0_184_29), .A1 (n_0_184_5), .A2 (n_0_184_14));
INV_X1 i_0_184_28 (.ZN (n_0_184_28), .A (n_0_184_14));
INV_X1 i_0_184_27 (.ZN (n_0_184_27), .A (n_0_184_5));
INV_X1 i_0_184_26 (.ZN (n_0_184_26), .A (n_0_184_25));
NAND2_X1 i_0_184_25 (.ZN (n_0_184_25), .A1 (n_0_184_10), .A2 (data[1]));
NAND2_X1 i_0_184_24 (.ZN (n_0_184_24), .A1 (n_0_184_30), .A2 (n_0_184_27));
NAND3_X1 i_0_184_23 (.ZN (n_0_184_23), .A1 (n_0_184_31), .A2 (n_0_184_28), .A3 (n_0_184_10));
INV_X1 i_0_184_22 (.ZN (n_0_184_22), .A (sps__n34));
INV_X1 i_0_184_21 (.ZN (n_0_184_21), .A (sps__n7));
INV_X1 i_0_184_20 (.ZN (n_0_184_20), .A (sps__n13));
INV_X1 i_0_184_19 (.ZN (n_0_184_19), .A (sps__n49));
NAND4_X1 i_0_184_18 (.ZN (n_0_184_18), .A1 (n_0_184_22), .A2 (n_0_184_21), .A3 (n_0_184_20), .A4 (n_0_184_19));
INV_X1 i_0_184_17 (.ZN (n_0_184_17), .A (sps__n61));
INV_X1 i_0_184_12 (.ZN (n_0_184_16), .A (sps__n73));
INV_X1 i_0_184_11 (.ZN (n_0_184_15), .A (sps__n85));
NAND4_X1 i_0_184_6 (.ZN (n_0_184_14), .A1 (n_0_184_17), .A2 (n_0_184_16), .A3 (n_0_184_15), .A4 (sps__n1));
INV_X1 i_0_184_5 (.ZN (n_0_184_13), .A (sps__n119));
INV_X1 i_0_184_4 (.ZN (n_0_184_12), .A (sps__n97));
NAND3_X1 i_0_184_1 (.ZN (n_0_184_11), .A1 (n_0_184_13), .A2 (n_0_184_12), .A3 (sps__n113));
INV_X1 i_0_184_0 (.ZN (n_0_184_10), .A (n_0_184_11));
INV_X1 i_0_184_16 (.ZN (n_0_184_9), .A (sps__n67));
INV_X1 i_0_184_15 (.ZN (n_0_184_8), .A (sps__n21));
INV_X1 i_0_184_14 (.ZN (n_0_184_7), .A (sps__n79));
INV_X1 i_0_184_13 (.ZN (n_0_184_6), .A (sps__n106));
NAND4_X1 i_0_184_3 (.ZN (n_0_184_5), .A1 (n_0_184_9), .A2 (n_0_184_8), .A3 (n_0_184_7), .A4 (n_0_184_6));
INV_X1 i_0_184_10 (.ZN (n_0_184_4), .A (sps__n57));
INV_X1 i_0_184_9 (.ZN (n_0_184_3), .A (sps__n27));
INV_X1 i_0_184_8 (.ZN (n_0_184_2), .A (sps__n44));
INV_X1 i_0_184_7 (.ZN (n_0_184_1), .A (sps__n93));
NAND4_X1 i_0_184_2 (.ZN (n_0_184_0), .A1 (n_0_184_4), .A2 (n_0_184_3), .A3 (n_0_184_2), .A4 (n_0_184_1));
NAND3_X1 i_0_167_36 (.ZN (n_0_181), .A1 (n_0_167_33), .A2 (n_0_167_34), .A3 (n_0_167_35));
NAND2_X1 i_0_167_35 (.ZN (n_0_167_35), .A1 (n_0_167_24), .A2 (\mem[4][1] ));
NAND2_X1 i_0_167_34 (.ZN (n_0_167_34), .A1 (n_0_167_23), .A2 (\mem[4][1] ));
NAND3_X1 i_0_167_33 (.ZN (n_0_167_33), .A1 (n_0_167_26), .A2 (n_0_167_32), .A3 (n_0_167_29));
NOR2_X1 i_0_167_32 (.ZN (n_0_167_32), .A1 (n_0_167_0), .A2 (n_0_167_18));
INV_X1 i_0_167_31 (.ZN (n_0_167_31), .A (n_0_167_18));
INV_X1 i_0_167_30 (.ZN (n_0_167_30), .A (n_0_167_0));
NOR2_X1 i_0_167_29 (.ZN (n_0_167_29), .A1 (n_0_167_5), .A2 (n_0_167_14));
INV_X1 i_0_167_28 (.ZN (n_0_167_28), .A (n_0_167_14));
INV_X1 i_0_167_27 (.ZN (n_0_167_27), .A (n_0_167_5));
INV_X1 i_0_167_26 (.ZN (n_0_167_26), .A (n_0_167_25));
NAND2_X1 i_0_167_25 (.ZN (n_0_167_25), .A1 (n_0_167_10), .A2 (data[1]));
NAND2_X1 i_0_167_24 (.ZN (n_0_167_24), .A1 (n_0_167_30), .A2 (n_0_167_27));
NAND3_X1 i_0_167_23 (.ZN (n_0_167_23), .A1 (n_0_167_31), .A2 (n_0_167_28), .A3 (n_0_167_10));
INV_X1 i_0_167_22 (.ZN (n_0_167_22), .A (sps__n34));
INV_X1 i_0_167_21 (.ZN (n_0_167_21), .A (sps__n7));
INV_X1 i_0_167_20 (.ZN (n_0_167_20), .A (sps__n13));
INV_X1 i_0_167_19 (.ZN (n_0_167_19), .A (sps__n49));
NAND4_X1 i_0_167_18 (.ZN (n_0_167_18), .A1 (n_0_167_22), .A2 (n_0_167_21), .A3 (n_0_167_20), .A4 (n_0_167_19));
INV_X1 i_0_167_17 (.ZN (n_0_167_17), .A (sps__n61));
INV_X1 i_0_167_12 (.ZN (n_0_167_16), .A (sps__n73));
INV_X1 i_0_167_11 (.ZN (n_0_167_15), .A (sps__n85));
NAND4_X1 i_0_167_6 (.ZN (n_0_167_14), .A1 (n_0_167_17), .A2 (n_0_167_16), .A3 (n_0_167_15), .A4 (sps__n1));
INV_X1 i_0_167_5 (.ZN (n_0_167_13), .A (sps__n113));
INV_X1 i_0_167_4 (.ZN (n_0_167_12), .A (address[0]));
NAND3_X1 i_0_167_1 (.ZN (n_0_167_11), .A1 (n_0_167_13), .A2 (n_0_167_12), .A3 (sps__n119));
INV_X1 i_0_167_0 (.ZN (n_0_167_10), .A (n_0_167_11));
INV_X1 i_0_167_16 (.ZN (n_0_167_9), .A (sps__n69));
INV_X1 i_0_167_15 (.ZN (n_0_167_8), .A (sps__n21));
INV_X1 i_0_167_14 (.ZN (n_0_167_7), .A (sps__n79));
INV_X1 i_0_167_13 (.ZN (n_0_167_6), .A (sps__n106));
NAND4_X1 i_0_167_3 (.ZN (n_0_167_5), .A1 (n_0_167_9), .A2 (n_0_167_8), .A3 (n_0_167_7), .A4 (n_0_167_6));
INV_X1 i_0_167_10 (.ZN (n_0_167_4), .A (sps__n56));
INV_X1 i_0_167_9 (.ZN (n_0_167_3), .A (sps__n27));
INV_X1 i_0_167_8 (.ZN (n_0_167_2), .A (sps__n41));
INV_X1 i_0_167_7 (.ZN (n_0_167_1), .A (sps__n93));
NAND4_X1 i_0_167_2 (.ZN (n_0_167_0), .A1 (n_0_167_4), .A2 (n_0_167_3), .A3 (n_0_167_2), .A4 (n_0_167_1));
NAND3_X1 i_0_133_35 (.ZN (n_0_180), .A1 (n_0_133_32), .A2 (n_0_133_33), .A3 (n_0_133_34));
NAND2_X1 i_0_133_34 (.ZN (n_0_133_34), .A1 (n_0_133_23), .A2 (\mem[8][2] ));
NAND3_X1 i_0_133_29 (.ZN (n_0_133_33), .A1 (n_0_133_26), .A2 (n_0_133_31), .A3 (n_0_133_28));
NAND2_X1 i_0_133_28 (.ZN (n_0_133_32), .A1 (n_0_133_27), .A2 (\mem[8][2] ));
NOR2_X1 i_0_133_24 (.ZN (n_0_133_31), .A1 (n_0_133_18), .A2 (n_0_133_0));
INV_X1 i_0_133_23 (.ZN (n_0_133_30), .A (n_0_133_0));
INV_X1 i_0_133_22 (.ZN (n_0_133_29), .A (n_0_133_18));
INV_X1 i_0_133_21 (.ZN (n_0_133_28), .A (n_0_133_5));
NAND3_X1 i_0_133_20 (.ZN (n_0_133_27), .A1 (n_0_133_28), .A2 (n_0_133_30), .A3 (n_0_133_9));
NOR2_X1 i_0_133_19 (.ZN (n_0_133_26), .A1 (n_0_133_14), .A2 (n_0_133_24));
INV_X1 i_0_133_18 (.ZN (n_0_133_25), .A (n_0_133_14));
NAND2_X1 i_0_133_17 (.ZN (n_0_133_24), .A1 (n_0_133_9), .A2 (data[2]));
NAND2_X1 i_0_133_16 (.ZN (n_0_133_23), .A1 (n_0_133_29), .A2 (n_0_133_25));
INV_X1 i_0_133_33 (.ZN (n_0_133_22), .A (sps__n35));
INV_X1 i_0_133_32 (.ZN (n_0_133_21), .A (sps__n8));
INV_X1 i_0_133_31 (.ZN (n_0_133_20), .A (sps__n13));
INV_X1 i_0_133_30 (.ZN (n_0_133_19), .A (sps__n50));
NAND4_X1 i_0_133_3 (.ZN (n_0_133_18), .A1 (n_0_133_22), .A2 (n_0_133_21), .A3 (n_0_133_20), .A4 (n_0_133_19));
INV_X1 i_0_133_27 (.ZN (n_0_133_17), .A (sps__n63));
INV_X1 i_0_133_26 (.ZN (n_0_133_16), .A (sps__n75));
INV_X1 i_0_133_25 (.ZN (n_0_133_15), .A (sps__n87));
NAND4_X1 i_0_133_8 (.ZN (n_0_133_14), .A1 (n_0_133_17), .A2 (n_0_133_16), .A3 (n_0_133_15), .A4 (sps__n1));
INV_X1 i_0_133_15 (.ZN (n_0_133_13), .A (sps__n121));
INV_X1 i_0_133_14 (.ZN (n_0_133_12), .A (sps__n112));
INV_X1 i_0_133_13 (.ZN (n_0_133_11), .A (sps__n97));
NAND3_X1 i_0_133_12 (.ZN (n_0_133_10), .A1 (n_0_133_13), .A2 (n_0_133_12), .A3 (n_0_133_11));
INV_X1 i_0_133_11 (.ZN (n_0_133_9), .A (n_0_133_10));
INV_X1 i_0_133_10 (.ZN (n_0_133_8), .A (sps__n67));
INV_X1 i_0_133_9 (.ZN (n_0_133_7), .A (sps__n21));
INV_X1 i_0_133_7 (.ZN (n_0_133_6), .A (sps__n80));
NAND4_X1 i_0_133_6 (.ZN (n_0_133_5), .A1 (n_0_133_8), .A2 (n_0_133_7), .A3 (n_0_133_6), .A4 (sps__n106));
INV_X1 i_0_133_5 (.ZN (n_0_133_4), .A (sps__n57));
INV_X1 i_0_133_4 (.ZN (n_0_133_3), .A (sps__n27));
INV_X1 i_0_133_2 (.ZN (n_0_133_2), .A (sps__n44));
INV_X1 i_0_133_1 (.ZN (n_0_133_1), .A (sps__n93));
NAND4_X1 i_0_133_0 (.ZN (n_0_133_0), .A1 (n_0_133_4), .A2 (n_0_133_3), .A3 (n_0_133_2), .A4 (n_0_133_1));
NAND3_X1 i_0_64_37 (.ZN (n_0_179), .A1 (n_0_64_34), .A2 (n_0_64_35), .A3 (n_0_64_36));
NAND2_X1 i_0_64_36 (.ZN (n_0_64_36), .A1 (n_0_64_25), .A2 (\mem[0][2] ));
NAND3_X1 i_0_64_35 (.ZN (n_0_64_35), .A1 (n_0_64_27), .A2 (n_0_64_33), .A3 (n_0_64_30));
NAND2_X1 i_0_64_34 (.ZN (n_0_64_34), .A1 (n_0_64_24), .A2 (\mem[0][2] ));
NOR2_X1 i_0_64_33 (.ZN (n_0_64_33), .A1 (n_0_64_0), .A2 (n_0_64_19));
INV_X1 i_0_64_32 (.ZN (n_0_64_32), .A (n_0_64_19));
INV_X1 i_0_64_31 (.ZN (n_0_64_31), .A (n_0_64_0));
NOR2_X1 i_0_64_30 (.ZN (n_0_64_30), .A1 (n_0_64_5), .A2 (n_0_64_15));
INV_X1 i_0_64_29 (.ZN (n_0_64_29), .A (n_0_64_15));
INV_X1 i_0_64_28 (.ZN (n_0_64_28), .A (n_0_64_5));
INV_X1 i_0_64_27 (.ZN (n_0_64_27), .A (n_0_64_26));
NAND2_X1 i_0_64_26 (.ZN (n_0_64_26), .A1 (n_0_64_10), .A2 (data[2]));
NAND2_X1 i_0_64_25 (.ZN (n_0_64_25), .A1 (n_0_64_31), .A2 (n_0_64_28));
NAND3_X1 i_0_64_24 (.ZN (n_0_64_24), .A1 (n_0_64_32), .A2 (n_0_64_29), .A3 (n_0_64_10));
INV_X1 i_0_64_23 (.ZN (n_0_64_23), .A (sps__n34));
INV_X1 i_0_64_22 (.ZN (n_0_64_22), .A (sps__n8));
INV_X1 i_0_64_21 (.ZN (n_0_64_21), .A (sps__n14));
INV_X1 i_0_64_20 (.ZN (n_0_64_20), .A (sps__n50));
NAND4_X1 i_0_64_19 (.ZN (n_0_64_19), .A1 (n_0_64_23), .A2 (n_0_64_22), .A3 (n_0_64_21), .A4 (n_0_64_20));
INV_X1 i_0_64_18 (.ZN (n_0_64_18), .A (sps__n63));
INV_X1 i_0_64_17 (.ZN (n_0_64_17), .A (sps__n75));
INV_X1 i_0_64_12 (.ZN (n_0_64_16), .A (sps__n87));
NAND4_X1 i_0_64_11 (.ZN (n_0_64_15), .A1 (n_0_64_18), .A2 (n_0_64_17), .A3 (n_0_64_16), .A4 (sps__n3));
INV_X1 i_0_64_6 (.ZN (n_0_64_14), .A (sps__n121));
INV_X1 i_0_64_5 (.ZN (n_0_64_13), .A (sps__n112));
INV_X1 i_0_64_4 (.ZN (n_0_64_12), .A (sps__n99));
NAND3_X1 i_0_64_1 (.ZN (n_0_64_11), .A1 (n_0_64_14), .A2 (n_0_64_13), .A3 (n_0_64_12));
INV_X1 i_0_64_0 (.ZN (n_0_64_10), .A (n_0_64_11));
INV_X1 i_0_64_16 (.ZN (n_0_64_9), .A (sps__n67));
INV_X1 i_0_64_15 (.ZN (n_0_64_8), .A (sps__n19));
INV_X1 i_0_64_14 (.ZN (n_0_64_7), .A (sps__n81));
INV_X1 i_0_64_13 (.ZN (n_0_64_6), .A (sps__n104));
NAND4_X1 i_0_64_3 (.ZN (n_0_64_5), .A1 (n_0_64_9), .A2 (n_0_64_8), .A3 (n_0_64_7), .A4 (n_0_64_6));
INV_X1 i_0_64_10 (.ZN (n_0_64_4), .A (sps__n57));
INV_X1 i_0_64_9 (.ZN (n_0_64_3), .A (sps__n26));
INV_X1 i_0_64_8 (.ZN (n_0_64_2), .A (sps__n43));
INV_X1 i_0_64_7 (.ZN (n_0_64_1), .A (sps__n91));
NAND4_X1 i_0_64_2 (.ZN (n_0_64_0), .A1 (n_0_64_4), .A2 (n_0_64_3), .A3 (n_0_64_2), .A4 (n_0_64_1));
NAND3_X1 i_0_198_37 (.ZN (n_0_178), .A1 (n_0_198_34), .A2 (n_0_198_35), .A3 (n_0_198_36));
NAND2_X1 i_0_198_36 (.ZN (n_0_198_36), .A1 (n_0_198_25), .A2 (\mem[0][3] ));
NAND3_X1 i_0_198_35 (.ZN (n_0_198_35), .A1 (n_0_198_27), .A2 (n_0_198_33), .A3 (n_0_198_30));
NAND2_X1 i_0_198_34 (.ZN (n_0_198_34), .A1 (n_0_198_24), .A2 (\mem[0][3] ));
NOR2_X1 i_0_198_33 (.ZN (n_0_198_33), .A1 (n_0_198_0), .A2 (n_0_198_19));
INV_X1 i_0_198_32 (.ZN (n_0_198_32), .A (n_0_198_19));
INV_X1 i_0_198_31 (.ZN (n_0_198_31), .A (n_0_198_0));
NOR2_X1 i_0_198_30 (.ZN (n_0_198_30), .A1 (n_0_198_5), .A2 (n_0_198_15));
INV_X1 i_0_198_29 (.ZN (n_0_198_29), .A (n_0_198_15));
INV_X1 i_0_198_28 (.ZN (n_0_198_28), .A (n_0_198_5));
INV_X1 i_0_198_27 (.ZN (n_0_198_27), .A (n_0_198_26));
NAND2_X1 i_0_198_26 (.ZN (n_0_198_26), .A1 (n_0_198_10), .A2 (data[3]));
NAND2_X1 i_0_198_25 (.ZN (n_0_198_25), .A1 (n_0_198_31), .A2 (n_0_198_28));
NAND3_X1 i_0_198_24 (.ZN (n_0_198_24), .A1 (n_0_198_32), .A2 (n_0_198_29), .A3 (n_0_198_10));
INV_X1 i_0_198_23 (.ZN (n_0_198_23), .A (sps__n34));
INV_X1 i_0_198_22 (.ZN (n_0_198_22), .A (sps__n9));
INV_X1 i_0_198_21 (.ZN (n_0_198_21), .A (sps__n15));
INV_X1 i_0_198_20 (.ZN (n_0_198_20), .A (sps__n51));
NAND4_X1 i_0_198_19 (.ZN (n_0_198_19), .A1 (n_0_198_23), .A2 (n_0_198_22), .A3 (n_0_198_21), .A4 (n_0_198_20));
INV_X1 i_0_198_18 (.ZN (n_0_198_18), .A (sps__n62));
INV_X1 i_0_198_17 (.ZN (n_0_198_17), .A (sps__n74));
INV_X1 i_0_198_12 (.ZN (n_0_198_16), .A (sps__n86));
NAND4_X1 i_0_198_11 (.ZN (n_0_198_15), .A1 (n_0_198_18), .A2 (n_0_198_17), .A3 (n_0_198_16), .A4 (sps__n3));
INV_X1 i_0_198_6 (.ZN (n_0_198_14), .A (sps__n122));
INV_X1 i_0_198_5 (.ZN (n_0_198_13), .A (sps__n112));
INV_X1 i_0_198_4 (.ZN (n_0_198_12), .A (sps__n99));
NAND3_X1 i_0_198_1 (.ZN (n_0_198_11), .A1 (n_0_198_14), .A2 (n_0_198_13), .A3 (n_0_198_12));
INV_X1 i_0_198_0 (.ZN (n_0_198_10), .A (n_0_198_11));
INV_X1 i_0_198_16 (.ZN (n_0_198_9), .A (sps__n67));
INV_X1 i_0_198_15 (.ZN (n_0_198_8), .A (sps__n19));
INV_X1 i_0_198_14 (.ZN (n_0_198_7), .A (sps__n81));
INV_X1 i_0_198_13 (.ZN (n_0_198_6), .A (sps__n105));
NAND4_X1 i_0_198_3 (.ZN (n_0_198_5), .A1 (n_0_198_9), .A2 (n_0_198_8), .A3 (n_0_198_7), .A4 (n_0_198_6));
INV_X1 i_0_198_10 (.ZN (n_0_198_4), .A (sps__n55));
INV_X1 i_0_198_9 (.ZN (n_0_198_3), .A (sps__n28));
INV_X1 i_0_198_8 (.ZN (n_0_198_2), .A (sps__n43));
INV_X1 i_0_198_7 (.ZN (n_0_198_1), .A (sps__n92));
NAND4_X1 i_0_198_2 (.ZN (n_0_198_0), .A1 (n_0_198_4), .A2 (n_0_198_3), .A3 (n_0_198_2), .A4 (n_0_198_1));
NAND3_X1 i_0_197_37 (.ZN (n_0_177), .A1 (n_0_197_34), .A2 (n_0_197_35), .A3 (n_0_197_36));
NAND2_X1 i_0_197_36 (.ZN (n_0_197_36), .A1 (n_0_197_25), .A2 (\mem[0][4] ));
NAND3_X1 i_0_197_35 (.ZN (n_0_197_35), .A1 (n_0_197_27), .A2 (n_0_197_33), .A3 (n_0_197_30));
NAND2_X1 i_0_197_34 (.ZN (n_0_197_34), .A1 (n_0_197_24), .A2 (\mem[0][4] ));
NOR2_X1 i_0_197_33 (.ZN (n_0_197_33), .A1 (n_0_197_0), .A2 (n_0_197_19));
INV_X1 i_0_197_32 (.ZN (n_0_197_32), .A (n_0_197_19));
INV_X1 i_0_197_31 (.ZN (n_0_197_31), .A (n_0_197_0));
NOR2_X1 i_0_197_30 (.ZN (n_0_197_30), .A1 (n_0_197_5), .A2 (n_0_197_15));
INV_X1 i_0_197_29 (.ZN (n_0_197_29), .A (n_0_197_15));
INV_X1 i_0_197_28 (.ZN (n_0_197_28), .A (n_0_197_5));
INV_X1 i_0_197_27 (.ZN (n_0_197_27), .A (n_0_197_26));
NAND2_X1 i_0_197_26 (.ZN (n_0_197_26), .A1 (n_0_197_10), .A2 (data[4]));
NAND2_X1 i_0_197_25 (.ZN (n_0_197_25), .A1 (n_0_197_31), .A2 (n_0_197_28));
NAND3_X1 i_0_197_24 (.ZN (n_0_197_24), .A1 (n_0_197_32), .A2 (n_0_197_29), .A3 (n_0_197_10));
INV_X1 i_0_197_23 (.ZN (n_0_197_23), .A (sps__n34));
INV_X1 i_0_197_22 (.ZN (n_0_197_22), .A (sps__n9));
INV_X1 i_0_197_21 (.ZN (n_0_197_21), .A (sps__n15));
INV_X1 i_0_197_20 (.ZN (n_0_197_20), .A (sps__n51));
NAND4_X1 i_0_197_19 (.ZN (n_0_197_19), .A1 (n_0_197_23), .A2 (n_0_197_22), .A3 (n_0_197_21), .A4 (n_0_197_20));
INV_X1 i_0_197_18 (.ZN (n_0_197_18), .A (sps__n62));
INV_X1 i_0_197_17 (.ZN (n_0_197_17), .A (sps__n75));
INV_X1 i_0_197_12 (.ZN (n_0_197_16), .A (sps__n86));
NAND4_X1 i_0_197_11 (.ZN (n_0_197_15), .A1 (n_0_197_18), .A2 (n_0_197_17), .A3 (n_0_197_16), .A4 (sps__n3));
INV_X1 i_0_197_6 (.ZN (n_0_197_14), .A (sps__n122));
INV_X1 i_0_197_5 (.ZN (n_0_197_13), .A (sps__n112));
INV_X1 i_0_197_4 (.ZN (n_0_197_12), .A (sps__n99));
NAND3_X1 i_0_197_1 (.ZN (n_0_197_11), .A1 (n_0_197_14), .A2 (n_0_197_13), .A3 (n_0_197_12));
INV_X1 i_0_197_0 (.ZN (n_0_197_10), .A (n_0_197_11));
INV_X1 i_0_197_16 (.ZN (n_0_197_9), .A (sps__n67));
INV_X1 i_0_197_15 (.ZN (n_0_197_8), .A (sps__n19));
INV_X1 i_0_197_14 (.ZN (n_0_197_7), .A (sps__n81));
INV_X1 i_0_197_13 (.ZN (n_0_197_6), .A (sps__n104));
NAND4_X1 i_0_197_3 (.ZN (n_0_197_5), .A1 (n_0_197_9), .A2 (n_0_197_8), .A3 (n_0_197_7), .A4 (n_0_197_6));
INV_X1 i_0_197_10 (.ZN (n_0_197_4), .A (sps__n55));
INV_X1 i_0_197_9 (.ZN (n_0_197_3), .A (sps__n28));
INV_X1 i_0_197_8 (.ZN (n_0_197_2), .A (sps__n43));
INV_X1 i_0_197_7 (.ZN (n_0_197_1), .A (sps__n92));
NAND4_X1 i_0_197_2 (.ZN (n_0_197_0), .A1 (n_0_197_4), .A2 (n_0_197_3), .A3 (n_0_197_2), .A4 (n_0_197_1));
NAND3_X1 i_0_169_36 (.ZN (n_0_176), .A1 (n_0_169_33), .A2 (n_0_169_34), .A3 (n_0_169_35));
NAND2_X1 i_0_169_35 (.ZN (n_0_169_35), .A1 (n_0_169_24), .A2 (\mem[1][2] ));
NAND2_X1 i_0_169_34 (.ZN (n_0_169_34), .A1 (n_0_169_23), .A2 (\mem[1][2] ));
NAND3_X1 i_0_169_33 (.ZN (n_0_169_33), .A1 (n_0_169_26), .A2 (n_0_169_32), .A3 (n_0_169_29));
NOR2_X1 i_0_169_32 (.ZN (n_0_169_32), .A1 (n_0_169_0), .A2 (n_0_169_18));
INV_X1 i_0_169_31 (.ZN (n_0_169_31), .A (n_0_169_18));
INV_X1 i_0_169_30 (.ZN (n_0_169_30), .A (n_0_169_0));
NOR2_X1 i_0_169_29 (.ZN (n_0_169_29), .A1 (n_0_169_5), .A2 (n_0_169_14));
INV_X1 i_0_169_28 (.ZN (n_0_169_28), .A (n_0_169_14));
INV_X1 i_0_169_27 (.ZN (n_0_169_27), .A (n_0_169_5));
INV_X1 i_0_169_26 (.ZN (n_0_169_26), .A (n_0_169_25));
NAND2_X1 i_0_169_25 (.ZN (n_0_169_25), .A1 (n_0_169_10), .A2 (data[2]));
NAND2_X1 i_0_169_24 (.ZN (n_0_169_24), .A1 (n_0_169_30), .A2 (n_0_169_27));
NAND3_X1 i_0_169_23 (.ZN (n_0_169_23), .A1 (n_0_169_31), .A2 (n_0_169_28), .A3 (n_0_169_10));
INV_X1 i_0_169_22 (.ZN (n_0_169_22), .A (sps__n34));
INV_X1 i_0_169_21 (.ZN (n_0_169_21), .A (sps__n8));
INV_X1 i_0_169_20 (.ZN (n_0_169_20), .A (sps__n14));
INV_X1 i_0_169_19 (.ZN (n_0_169_19), .A (sps__n50));
NAND4_X1 i_0_169_18 (.ZN (n_0_169_18), .A1 (n_0_169_22), .A2 (n_0_169_21), .A3 (n_0_169_20), .A4 (n_0_169_19));
INV_X1 i_0_169_17 (.ZN (n_0_169_17), .A (sps__n63));
INV_X1 i_0_169_12 (.ZN (n_0_169_16), .A (sps__n74));
INV_X1 i_0_169_11 (.ZN (n_0_169_15), .A (sps__n87));
NAND4_X1 i_0_169_6 (.ZN (n_0_169_14), .A1 (n_0_169_17), .A2 (n_0_169_16), .A3 (n_0_169_15), .A4 (sps__n3));
INV_X1 i_0_169_5 (.ZN (n_0_169_13), .A (sps__n121));
INV_X1 i_0_169_4 (.ZN (n_0_169_12), .A (sps__n112));
NAND3_X1 i_0_169_1 (.ZN (n_0_169_11), .A1 (n_0_169_13), .A2 (n_0_169_12), .A3 (sps__n99));
INV_X1 i_0_169_0 (.ZN (n_0_169_10), .A (n_0_169_11));
INV_X1 i_0_169_16 (.ZN (n_0_169_9), .A (sps__n67));
INV_X1 i_0_169_15 (.ZN (n_0_169_8), .A (sps__n19));
INV_X1 i_0_169_14 (.ZN (n_0_169_7), .A (sps__n81));
INV_X1 i_0_169_13 (.ZN (n_0_169_6), .A (sps__n104));
NAND4_X1 i_0_169_3 (.ZN (n_0_169_5), .A1 (n_0_169_9), .A2 (n_0_169_8), .A3 (n_0_169_7), .A4 (n_0_169_6));
INV_X1 i_0_169_10 (.ZN (n_0_169_4), .A (sps__n57));
INV_X1 i_0_169_9 (.ZN (n_0_169_3), .A (sps__n26));
INV_X1 i_0_169_8 (.ZN (n_0_169_2), .A (sps__n43));
INV_X1 i_0_169_7 (.ZN (n_0_169_1), .A (sps__n91));
NAND4_X1 i_0_169_2 (.ZN (n_0_169_0), .A1 (n_0_169_4), .A2 (n_0_169_3), .A3 (n_0_169_2), .A4 (n_0_169_1));
NAND3_X1 i_0_183_36 (.ZN (n_0_175), .A1 (n_0_183_33), .A2 (n_0_183_34), .A3 (n_0_183_35));
NAND2_X1 i_0_183_35 (.ZN (n_0_183_35), .A1 (n_0_183_24), .A2 (\mem[1][3] ));
NAND2_X1 i_0_183_34 (.ZN (n_0_183_34), .A1 (n_0_183_23), .A2 (\mem[1][3] ));
NAND3_X1 i_0_183_33 (.ZN (n_0_183_33), .A1 (n_0_183_26), .A2 (n_0_183_32), .A3 (n_0_183_29));
NOR2_X1 i_0_183_32 (.ZN (n_0_183_32), .A1 (n_0_183_0), .A2 (n_0_183_18));
INV_X1 i_0_183_31 (.ZN (n_0_183_31), .A (n_0_183_18));
INV_X1 i_0_183_30 (.ZN (n_0_183_30), .A (n_0_183_0));
NOR2_X1 i_0_183_29 (.ZN (n_0_183_29), .A1 (n_0_183_5), .A2 (n_0_183_14));
INV_X1 i_0_183_28 (.ZN (n_0_183_28), .A (n_0_183_14));
INV_X1 i_0_183_27 (.ZN (n_0_183_27), .A (n_0_183_5));
INV_X1 i_0_183_26 (.ZN (n_0_183_26), .A (n_0_183_25));
NAND2_X1 i_0_183_25 (.ZN (n_0_183_25), .A1 (n_0_183_10), .A2 (data[3]));
NAND2_X1 i_0_183_24 (.ZN (n_0_183_24), .A1 (n_0_183_30), .A2 (n_0_183_27));
NAND3_X1 i_0_183_23 (.ZN (n_0_183_23), .A1 (n_0_183_31), .A2 (n_0_183_28), .A3 (n_0_183_10));
INV_X1 i_0_183_22 (.ZN (n_0_183_22), .A (sps__n34));
INV_X1 i_0_183_21 (.ZN (n_0_183_21), .A (sps__n8));
INV_X1 i_0_183_20 (.ZN (n_0_183_20), .A (sps__n14));
INV_X1 i_0_183_19 (.ZN (n_0_183_19), .A (sps__n50));
NAND4_X1 i_0_183_18 (.ZN (n_0_183_18), .A1 (n_0_183_22), .A2 (n_0_183_21), .A3 (n_0_183_20), .A4 (n_0_183_19));
INV_X1 i_0_183_17 (.ZN (n_0_183_17), .A (sps__n63));
INV_X1 i_0_183_12 (.ZN (n_0_183_16), .A (sps__n74));
INV_X1 i_0_183_11 (.ZN (n_0_183_15), .A (sps__n87));
NAND4_X1 i_0_183_6 (.ZN (n_0_183_14), .A1 (n_0_183_17), .A2 (n_0_183_16), .A3 (n_0_183_15), .A4 (sps__n3));
INV_X1 i_0_183_5 (.ZN (n_0_183_13), .A (sps__n121));
INV_X1 i_0_183_4 (.ZN (n_0_183_12), .A (sps__n112));
NAND3_X1 i_0_183_1 (.ZN (n_0_183_11), .A1 (n_0_183_13), .A2 (n_0_183_12), .A3 (sps__n99));
INV_X1 i_0_183_0 (.ZN (n_0_183_10), .A (n_0_183_11));
INV_X1 i_0_183_16 (.ZN (n_0_183_9), .A (sps__n68));
INV_X1 i_0_183_15 (.ZN (n_0_183_8), .A (sps__n21));
INV_X1 i_0_183_14 (.ZN (n_0_183_7), .A (sps__n80));
INV_X1 i_0_183_13 (.ZN (n_0_183_6), .A (sps__n103));
NAND4_X1 i_0_183_3 (.ZN (n_0_183_5), .A1 (n_0_183_9), .A2 (n_0_183_8), .A3 (n_0_183_7), .A4 (n_0_183_6));
INV_X1 i_0_183_10 (.ZN (n_0_183_4), .A (sps__n57));
INV_X1 i_0_183_9 (.ZN (n_0_183_3), .A (sps__n26));
INV_X1 i_0_183_8 (.ZN (n_0_183_2), .A (sps__n44));
INV_X1 i_0_183_7 (.ZN (n_0_183_1), .A (sps__n91));
NAND4_X1 i_0_183_2 (.ZN (n_0_183_0), .A1 (n_0_183_4), .A2 (n_0_183_3), .A3 (n_0_183_2), .A4 (n_0_183_1));
NAND3_X1 i_0_182_36 (.ZN (n_0_174), .A1 (n_0_182_33), .A2 (n_0_182_34), .A3 (n_0_182_35));
NAND2_X1 i_0_182_35 (.ZN (n_0_182_35), .A1 (n_0_182_24), .A2 (\mem[1][4] ));
NAND2_X1 i_0_182_34 (.ZN (n_0_182_34), .A1 (n_0_182_23), .A2 (\mem[1][4] ));
NAND3_X1 i_0_182_33 (.ZN (n_0_182_33), .A1 (n_0_182_26), .A2 (n_0_182_32), .A3 (n_0_182_29));
NOR2_X1 i_0_182_32 (.ZN (n_0_182_32), .A1 (n_0_182_0), .A2 (n_0_182_18));
INV_X1 i_0_182_31 (.ZN (n_0_182_31), .A (n_0_182_18));
INV_X1 i_0_182_30 (.ZN (n_0_182_30), .A (n_0_182_0));
NOR2_X1 i_0_182_29 (.ZN (n_0_182_29), .A1 (n_0_182_5), .A2 (n_0_182_14));
INV_X1 i_0_182_28 (.ZN (n_0_182_28), .A (n_0_182_14));
INV_X1 i_0_182_27 (.ZN (n_0_182_27), .A (n_0_182_5));
INV_X1 i_0_182_26 (.ZN (n_0_182_26), .A (n_0_182_25));
NAND2_X1 i_0_182_25 (.ZN (n_0_182_25), .A1 (n_0_182_10), .A2 (data[4]));
NAND2_X1 i_0_182_24 (.ZN (n_0_182_24), .A1 (n_0_182_30), .A2 (n_0_182_27));
NAND3_X1 i_0_182_23 (.ZN (n_0_182_23), .A1 (n_0_182_31), .A2 (n_0_182_28), .A3 (n_0_182_10));
INV_X1 i_0_182_22 (.ZN (n_0_182_22), .A (sps__n34));
INV_X1 i_0_182_21 (.ZN (n_0_182_21), .A (sps__n8));
INV_X1 i_0_182_20 (.ZN (n_0_182_20), .A (sps__n14));
INV_X1 i_0_182_19 (.ZN (n_0_182_19), .A (sps__n50));
NAND4_X1 i_0_182_18 (.ZN (n_0_182_18), .A1 (n_0_182_22), .A2 (n_0_182_21), .A3 (n_0_182_20), .A4 (n_0_182_19));
INV_X1 i_0_182_17 (.ZN (n_0_182_17), .A (sps__n63));
INV_X1 i_0_182_12 (.ZN (n_0_182_16), .A (sps__n74));
INV_X1 i_0_182_11 (.ZN (n_0_182_15), .A (sps__n87));
NAND4_X1 i_0_182_6 (.ZN (n_0_182_14), .A1 (n_0_182_17), .A2 (n_0_182_16), .A3 (n_0_182_15), .A4 (sps__n3));
INV_X1 i_0_182_5 (.ZN (n_0_182_13), .A (sps__n122));
INV_X1 i_0_182_4 (.ZN (n_0_182_12), .A (sps__n112));
NAND3_X1 i_0_182_1 (.ZN (n_0_182_11), .A1 (n_0_182_13), .A2 (n_0_182_12), .A3 (sps__n99));
INV_X1 i_0_182_0 (.ZN (n_0_182_10), .A (n_0_182_11));
INV_X1 i_0_182_16 (.ZN (n_0_182_9), .A (sps__n67));
INV_X1 i_0_182_15 (.ZN (n_0_182_8), .A (sps__n19));
INV_X1 i_0_182_14 (.ZN (n_0_182_7), .A (sps__n81));
INV_X1 i_0_182_13 (.ZN (n_0_182_6), .A (sps__n104));
NAND4_X1 i_0_182_3 (.ZN (n_0_182_5), .A1 (n_0_182_9), .A2 (n_0_182_8), .A3 (n_0_182_7), .A4 (n_0_182_6));
INV_X1 i_0_182_10 (.ZN (n_0_182_4), .A (sps__n57));
INV_X1 i_0_182_9 (.ZN (n_0_182_3), .A (sps__n26));
INV_X1 i_0_182_8 (.ZN (n_0_182_2), .A (sps__n43));
INV_X1 i_0_182_7 (.ZN (n_0_182_1), .A (sps__n91));
NAND4_X1 i_0_182_2 (.ZN (n_0_182_0), .A1 (n_0_182_4), .A2 (n_0_182_3), .A3 (n_0_182_2), .A4 (n_0_182_1));
NAND3_X1 i_0_181_36 (.ZN (n_0_173), .A1 (n_0_181_33), .A2 (n_0_181_34), .A3 (n_0_181_35));
NAND2_X1 i_0_181_35 (.ZN (n_0_181_35), .A1 (n_0_181_24), .A2 (\mem[2][2] ));
NAND2_X1 i_0_181_34 (.ZN (n_0_181_34), .A1 (n_0_181_23), .A2 (\mem[2][2] ));
NAND3_X1 i_0_181_33 (.ZN (n_0_181_33), .A1 (n_0_181_26), .A2 (n_0_181_32), .A3 (n_0_181_29));
NOR2_X1 i_0_181_32 (.ZN (n_0_181_32), .A1 (n_0_181_0), .A2 (n_0_181_18));
INV_X1 i_0_181_31 (.ZN (n_0_181_31), .A (n_0_181_18));
INV_X1 i_0_181_30 (.ZN (n_0_181_30), .A (n_0_181_0));
NOR2_X1 i_0_181_29 (.ZN (n_0_181_29), .A1 (n_0_181_5), .A2 (n_0_181_14));
INV_X1 i_0_181_28 (.ZN (n_0_181_28), .A (n_0_181_14));
INV_X1 i_0_181_27 (.ZN (n_0_181_27), .A (n_0_181_5));
INV_X1 i_0_181_26 (.ZN (n_0_181_26), .A (n_0_181_25));
NAND2_X1 i_0_181_25 (.ZN (n_0_181_25), .A1 (n_0_181_10), .A2 (data[2]));
NAND2_X1 i_0_181_24 (.ZN (n_0_181_24), .A1 (n_0_181_30), .A2 (n_0_181_27));
NAND3_X1 i_0_181_23 (.ZN (n_0_181_23), .A1 (n_0_181_31), .A2 (n_0_181_28), .A3 (n_0_181_10));
INV_X1 i_0_181_22 (.ZN (n_0_181_22), .A (sps__n35));
INV_X1 i_0_181_21 (.ZN (n_0_181_21), .A (sps__n8));
INV_X1 i_0_181_20 (.ZN (n_0_181_20), .A (sps__n13));
INV_X1 i_0_181_19 (.ZN (n_0_181_19), .A (sps__n50));
NAND4_X1 i_0_181_18 (.ZN (n_0_181_18), .A1 (n_0_181_22), .A2 (n_0_181_21), .A3 (n_0_181_20), .A4 (n_0_181_19));
INV_X1 i_0_181_17 (.ZN (n_0_181_17), .A (sps__n63));
INV_X1 i_0_181_12 (.ZN (n_0_181_16), .A (sps__n75));
INV_X1 i_0_181_11 (.ZN (n_0_181_15), .A (sps__n87));
NAND4_X1 i_0_181_6 (.ZN (n_0_181_14), .A1 (n_0_181_17), .A2 (n_0_181_16), .A3 (n_0_181_15), .A4 (sps__n1));
INV_X1 i_0_181_5 (.ZN (n_0_181_13), .A (sps__n121));
INV_X1 i_0_181_4 (.ZN (n_0_181_12), .A (sps__n97));
NAND3_X1 i_0_181_1 (.ZN (n_0_181_11), .A1 (n_0_181_13), .A2 (n_0_181_12), .A3 (sps__n112));
INV_X1 i_0_181_0 (.ZN (n_0_181_10), .A (n_0_181_11));
INV_X1 i_0_181_16 (.ZN (n_0_181_9), .A (sps__n67));
INV_X1 i_0_181_15 (.ZN (n_0_181_8), .A (sps__n21));
INV_X1 i_0_181_14 (.ZN (n_0_181_7), .A (sps__n80));
INV_X1 i_0_181_13 (.ZN (n_0_181_6), .A (sps__n103));
NAND4_X1 i_0_181_3 (.ZN (n_0_181_5), .A1 (n_0_181_9), .A2 (n_0_181_8), .A3 (n_0_181_7), .A4 (n_0_181_6));
INV_X1 i_0_181_10 (.ZN (n_0_181_4), .A (sps__n57));
INV_X1 i_0_181_9 (.ZN (n_0_181_3), .A (sps__n27));
INV_X1 i_0_181_8 (.ZN (n_0_181_2), .A (sps__n44));
INV_X1 i_0_181_7 (.ZN (n_0_181_1), .A (sps__n91));
NAND4_X1 i_0_181_2 (.ZN (n_0_181_0), .A1 (n_0_181_4), .A2 (n_0_181_3), .A3 (n_0_181_2), .A4 (n_0_181_1));
NAND3_X1 i_0_166_36 (.ZN (n_0_172), .A1 (n_0_166_33), .A2 (n_0_166_34), .A3 (n_0_166_35));
NAND2_X1 i_0_166_35 (.ZN (n_0_166_35), .A1 (n_0_166_24), .A2 (\mem[2][3] ));
NAND2_X1 i_0_166_34 (.ZN (n_0_166_34), .A1 (n_0_166_23), .A2 (\mem[2][3] ));
NAND3_X1 i_0_166_33 (.ZN (n_0_166_33), .A1 (n_0_166_26), .A2 (n_0_166_32), .A3 (n_0_166_29));
NOR2_X1 i_0_166_32 (.ZN (n_0_166_32), .A1 (n_0_166_0), .A2 (n_0_166_18));
INV_X1 i_0_166_31 (.ZN (n_0_166_31), .A (n_0_166_18));
INV_X1 i_0_166_30 (.ZN (n_0_166_30), .A (n_0_166_0));
NOR2_X1 i_0_166_29 (.ZN (n_0_166_29), .A1 (n_0_166_5), .A2 (n_0_166_14));
INV_X1 i_0_166_28 (.ZN (n_0_166_28), .A (n_0_166_14));
INV_X1 i_0_166_27 (.ZN (n_0_166_27), .A (n_0_166_5));
INV_X1 i_0_166_26 (.ZN (n_0_166_26), .A (n_0_166_25));
NAND2_X1 i_0_166_25 (.ZN (n_0_166_25), .A1 (n_0_166_10), .A2 (data[3]));
NAND2_X1 i_0_166_24 (.ZN (n_0_166_24), .A1 (n_0_166_30), .A2 (n_0_166_27));
NAND3_X1 i_0_166_23 (.ZN (n_0_166_23), .A1 (n_0_166_31), .A2 (n_0_166_28), .A3 (n_0_166_10));
INV_X1 i_0_166_22 (.ZN (n_0_166_22), .A (sps__n34));
INV_X1 i_0_166_21 (.ZN (n_0_166_21), .A (sps__n8));
INV_X1 i_0_166_20 (.ZN (n_0_166_20), .A (sps__n14));
INV_X1 i_0_166_19 (.ZN (n_0_166_19), .A (sps__n50));
NAND4_X1 i_0_166_18 (.ZN (n_0_166_18), .A1 (n_0_166_22), .A2 (n_0_166_21), .A3 (n_0_166_20), .A4 (n_0_166_19));
INV_X1 i_0_166_17 (.ZN (n_0_166_17), .A (sps__n63));
INV_X1 i_0_166_12 (.ZN (n_0_166_16), .A (sps__n74));
INV_X1 i_0_166_11 (.ZN (n_0_166_15), .A (sps__n86));
NAND4_X1 i_0_166_6 (.ZN (n_0_166_14), .A1 (n_0_166_17), .A2 (n_0_166_16), .A3 (n_0_166_15), .A4 (sps__n3));
INV_X1 i_0_166_5 (.ZN (n_0_166_13), .A (sps__n122));
INV_X1 i_0_166_4 (.ZN (n_0_166_12), .A (sps__n99));
NAND3_X1 i_0_166_1 (.ZN (n_0_166_11), .A1 (n_0_166_13), .A2 (n_0_166_12), .A3 (sps__n112));
INV_X1 i_0_166_0 (.ZN (n_0_166_10), .A (n_0_166_11));
INV_X1 i_0_166_16 (.ZN (n_0_166_9), .A (sps__n68));
INV_X1 i_0_166_15 (.ZN (n_0_166_8), .A (sps__n19));
INV_X1 i_0_166_14 (.ZN (n_0_166_7), .A (sps__n81));
INV_X1 i_0_166_13 (.ZN (n_0_166_6), .A (sps__n104));
NAND4_X1 i_0_166_3 (.ZN (n_0_166_5), .A1 (n_0_166_9), .A2 (n_0_166_8), .A3 (n_0_166_7), .A4 (n_0_166_6));
INV_X1 i_0_166_10 (.ZN (n_0_166_4), .A (sps__n57));
INV_X1 i_0_166_9 (.ZN (n_0_166_3), .A (sps__n26));
INV_X1 i_0_166_8 (.ZN (n_0_166_2), .A (sps__n43));
INV_X1 i_0_166_7 (.ZN (n_0_166_1), .A (sps__n91));
NAND4_X1 i_0_166_2 (.ZN (n_0_166_0), .A1 (n_0_166_4), .A2 (n_0_166_3), .A3 (n_0_166_2), .A4 (n_0_166_1));
NAND3_X1 i_0_165_36 (.ZN (n_0_171), .A1 (n_0_165_33), .A2 (n_0_165_34), .A3 (n_0_165_35));
NAND2_X1 i_0_165_35 (.ZN (n_0_165_35), .A1 (n_0_165_24), .A2 (\mem[2][4] ));
NAND2_X1 i_0_165_34 (.ZN (n_0_165_34), .A1 (n_0_165_23), .A2 (\mem[2][4] ));
NAND3_X1 i_0_165_33 (.ZN (n_0_165_33), .A1 (n_0_165_26), .A2 (n_0_165_32), .A3 (n_0_165_29));
NOR2_X1 i_0_165_32 (.ZN (n_0_165_32), .A1 (n_0_165_0), .A2 (n_0_165_18));
INV_X1 i_0_165_31 (.ZN (n_0_165_31), .A (n_0_165_18));
INV_X1 i_0_165_30 (.ZN (n_0_165_30), .A (n_0_165_0));
NOR2_X1 i_0_165_29 (.ZN (n_0_165_29), .A1 (n_0_165_5), .A2 (n_0_165_14));
INV_X1 i_0_165_28 (.ZN (n_0_165_28), .A (n_0_165_14));
INV_X1 i_0_165_27 (.ZN (n_0_165_27), .A (n_0_165_5));
INV_X1 i_0_165_26 (.ZN (n_0_165_26), .A (n_0_165_25));
NAND2_X1 i_0_165_25 (.ZN (n_0_165_25), .A1 (n_0_165_10), .A2 (data[4]));
NAND2_X1 i_0_165_24 (.ZN (n_0_165_24), .A1 (n_0_165_30), .A2 (n_0_165_27));
NAND3_X1 i_0_165_23 (.ZN (n_0_165_23), .A1 (n_0_165_31), .A2 (n_0_165_28), .A3 (n_0_165_10));
INV_X1 i_0_165_22 (.ZN (n_0_165_22), .A (sps__n34));
INV_X1 i_0_165_21 (.ZN (n_0_165_21), .A (sps__n8));
INV_X1 i_0_165_20 (.ZN (n_0_165_20), .A (sps__n14));
INV_X1 i_0_165_19 (.ZN (n_0_165_19), .A (sps__n50));
NAND4_X1 i_0_165_18 (.ZN (n_0_165_18), .A1 (n_0_165_22), .A2 (n_0_165_21), .A3 (n_0_165_20), .A4 (n_0_165_19));
INV_X1 i_0_165_17 (.ZN (n_0_165_17), .A (sps__n63));
INV_X1 i_0_165_12 (.ZN (n_0_165_16), .A (sps__n74));
INV_X1 i_0_165_11 (.ZN (n_0_165_15), .A (sps__n86));
NAND4_X1 i_0_165_6 (.ZN (n_0_165_14), .A1 (n_0_165_17), .A2 (n_0_165_16), .A3 (n_0_165_15), .A4 (sps__n3));
INV_X1 i_0_165_5 (.ZN (n_0_165_13), .A (sps__n122));
INV_X1 i_0_165_4 (.ZN (n_0_165_12), .A (sps__n99));
NAND3_X1 i_0_165_1 (.ZN (n_0_165_11), .A1 (n_0_165_13), .A2 (n_0_165_12), .A3 (sps__n112));
INV_X1 i_0_165_0 (.ZN (n_0_165_10), .A (n_0_165_11));
INV_X1 i_0_165_16 (.ZN (n_0_165_9), .A (sps__n67));
INV_X1 i_0_165_15 (.ZN (n_0_165_8), .A (sps__n19));
INV_X1 i_0_165_14 (.ZN (n_0_165_7), .A (sps__n81));
INV_X1 i_0_165_13 (.ZN (n_0_165_6), .A (sps__n104));
NAND4_X1 i_0_165_3 (.ZN (n_0_165_5), .A1 (n_0_165_9), .A2 (n_0_165_8), .A3 (n_0_165_7), .A4 (n_0_165_6));
INV_X1 i_0_165_10 (.ZN (n_0_165_4), .A (sps__n57));
INV_X1 i_0_165_9 (.ZN (n_0_165_3), .A (sps__n28));
INV_X1 i_0_165_8 (.ZN (n_0_165_2), .A (sps__n43));
INV_X1 i_0_165_7 (.ZN (n_0_165_1), .A (sps__n91));
NAND4_X1 i_0_165_2 (.ZN (n_0_165_0), .A1 (n_0_165_4), .A2 (n_0_165_3), .A3 (n_0_165_2), .A4 (n_0_165_1));
NAND3_X1 i_0_164_31 (.ZN (n_0_164_30), .A1 (n_0_164_27), .A2 (n_0_164_28), .A3 (n_0_164_29));
NOR2_X1 i_0_164_30 (.ZN (n_0_164_29), .A1 (n_0_164_13), .A2 (n_0_164_23));
NOR2_X1 i_0_164_29 (.ZN (n_0_164_28), .A1 (n_0_164_22), .A2 (n_0_164_21));
NOR2_X1 i_0_164_28 (.ZN (n_0_164_27), .A1 (n_0_164_17), .A2 (n_0_164_20));
NOR2_X1 i_0_164_27 (.ZN (n_0_164_26), .A1 (n_0_164_17), .A2 (n_0_164_13));
NOR2_X1 i_0_164_26 (.ZN (n_0_164_25), .A1 (n_0_164_20), .A2 (n_0_164_21));
NOR2_X1 i_0_164_25 (.ZN (n_0_164_24), .A1 (n_0_164_22), .A2 (n_0_164_23));
NAND3_X1 i_0_164_24 (.ZN (n_0_164_23), .A1 (n_0_164_4), .A2 (n_0_164_2), .A3 (n_0_164_6));
NAND3_X1 i_0_164_23 (.ZN (n_0_164_22), .A1 (n_0_164_1), .A2 (n_0_164_3), .A3 (n_0_164_5));
NAND3_X1 i_0_164_22 (.ZN (n_0_164_21), .A1 (n_0_164_10), .A2 (n_0_164_8), .A3 (n_0_164_12));
NAND3_X1 i_0_164_21 (.ZN (n_0_164_20), .A1 (n_0_164_7), .A2 (n_0_164_9), .A3 (n_0_164_11));
NAND2_X1 i_0_164_20 (.ZN (n_0_164_19), .A1 (n_0_164_30), .A2 (\mem[3][4] ));
INV_X1 i_0_164_19 (.ZN (n_0_164_18), .A (sps__n121));
NAND4_X1 i_0_164_18 (.ZN (n_0_164_17), .A1 (n_0_164_18), .A2 (sps__n1), .A3 (sps__n114), .A4 (sps__n97));
INV_X1 i_0_164_17 (.ZN (n_0_164_16), .A (sps__n21));
INV_X1 i_0_164_16 (.ZN (n_0_164_15), .A (sps__n80));
INV_X1 i_0_164_15 (.ZN (n_0_164_14), .A (sps__n103));
NAND3_X1 i_0_164_14 (.ZN (n_0_164_13), .A1 (n_0_164_16), .A2 (n_0_164_15), .A3 (n_0_164_14));
INV_X1 i_0_164_13 (.ZN (n_0_164_12), .A (sps__n61));
INV_X1 i_0_164_12 (.ZN (n_0_164_11), .A (sps__n74));
INV_X1 i_0_164_11 (.ZN (n_0_164_10), .A (sps__n7));
INV_X1 i_0_164_10 (.ZN (n_0_164_9), .A (sps__n13));
INV_X1 i_0_164_9 (.ZN (n_0_164_8), .A (sps__n87));
INV_X1 i_0_164_8 (.ZN (n_0_164_7), .A (sps__n36));
INV_X1 i_0_164_7 (.ZN (n_0_164_6), .A (sps__n91));
INV_X1 i_0_164_6 (.ZN (n_0_164_5), .A (sps__n69));
INV_X1 i_0_164_5 (.ZN (n_0_164_4), .A (sps__n27));
INV_X1 i_0_164_4 (.ZN (n_0_164_3), .A (sps__n41));
INV_X1 i_0_164_3 (.ZN (n_0_164_2), .A (sps__n49));
INV_X1 i_0_164_2 (.ZN (n_0_164_1), .A (sps__n56));
NAND4_X1 i_0_164_1 (.ZN (n_0_164_0), .A1 (n_0_164_26), .A2 (n_0_164_25), .A3 (n_0_164_24), .A4 (data[4]));
NAND2_X1 i_0_164_0 (.ZN (n_0_170), .A1 (n_0_164_19), .A2 (n_0_164_0));
NAND3_X1 i_0_147_36 (.ZN (n_0_169), .A1 (n_0_147_33), .A2 (n_0_147_34), .A3 (n_0_147_35));
NAND2_X1 i_0_147_35 (.ZN (n_0_147_35), .A1 (n_0_147_24), .A2 (\mem[4][2] ));
NAND2_X1 i_0_147_34 (.ZN (n_0_147_34), .A1 (n_0_147_23), .A2 (\mem[4][2] ));
NAND3_X1 i_0_147_33 (.ZN (n_0_147_33), .A1 (n_0_147_26), .A2 (n_0_147_32), .A3 (n_0_147_29));
NOR2_X1 i_0_147_32 (.ZN (n_0_147_32), .A1 (n_0_147_0), .A2 (n_0_147_18));
INV_X1 i_0_147_31 (.ZN (n_0_147_31), .A (n_0_147_18));
INV_X1 i_0_147_30 (.ZN (n_0_147_30), .A (n_0_147_0));
NOR2_X1 i_0_147_29 (.ZN (n_0_147_29), .A1 (n_0_147_5), .A2 (n_0_147_14));
INV_X1 i_0_147_28 (.ZN (n_0_147_28), .A (n_0_147_14));
INV_X1 i_0_147_27 (.ZN (n_0_147_27), .A (n_0_147_5));
INV_X1 i_0_147_26 (.ZN (n_0_147_26), .A (n_0_147_25));
NAND2_X1 i_0_147_25 (.ZN (n_0_147_25), .A1 (n_0_147_10), .A2 (data[2]));
NAND2_X1 i_0_147_24 (.ZN (n_0_147_24), .A1 (n_0_147_30), .A2 (n_0_147_27));
NAND3_X1 i_0_147_23 (.ZN (n_0_147_23), .A1 (n_0_147_31), .A2 (n_0_147_28), .A3 (n_0_147_10));
INV_X1 i_0_147_22 (.ZN (n_0_147_22), .A (sps__n34));
INV_X1 i_0_147_21 (.ZN (n_0_147_21), .A (sps__n8));
INV_X1 i_0_147_20 (.ZN (n_0_147_20), .A (sps__n14));
INV_X1 i_0_147_19 (.ZN (n_0_147_19), .A (sps__n50));
NAND4_X1 i_0_147_18 (.ZN (n_0_147_18), .A1 (n_0_147_22), .A2 (n_0_147_21), .A3 (n_0_147_20), .A4 (n_0_147_19));
INV_X1 i_0_147_17 (.ZN (n_0_147_17), .A (sps__n63));
INV_X1 i_0_147_12 (.ZN (n_0_147_16), .A (sps__n75));
INV_X1 i_0_147_11 (.ZN (n_0_147_15), .A (sps__n87));
NAND4_X1 i_0_147_6 (.ZN (n_0_147_14), .A1 (n_0_147_17), .A2 (n_0_147_16), .A3 (n_0_147_15), .A4 (sps__n3));
INV_X1 i_0_147_5 (.ZN (n_0_147_13), .A (sps__n112));
INV_X1 i_0_147_4 (.ZN (n_0_147_12), .A (sps__n99));
NAND3_X1 i_0_147_1 (.ZN (n_0_147_11), .A1 (n_0_147_13), .A2 (n_0_147_12), .A3 (sps__n121));
INV_X1 i_0_147_0 (.ZN (n_0_147_10), .A (n_0_147_11));
INV_X1 i_0_147_16 (.ZN (n_0_147_9), .A (sps__n67));
INV_X1 i_0_147_15 (.ZN (n_0_147_8), .A (sps__n19));
INV_X1 i_0_147_14 (.ZN (n_0_147_7), .A (sps__n81));
INV_X1 i_0_147_13 (.ZN (n_0_147_6), .A (sps__n104));
NAND4_X1 i_0_147_3 (.ZN (n_0_147_5), .A1 (n_0_147_9), .A2 (n_0_147_8), .A3 (n_0_147_7), .A4 (n_0_147_6));
INV_X1 i_0_147_10 (.ZN (n_0_147_4), .A (sps__n57));
INV_X1 i_0_147_9 (.ZN (n_0_147_3), .A (sps__n26));
INV_X1 i_0_147_8 (.ZN (n_0_147_2), .A (sps__n43));
INV_X1 i_0_147_7 (.ZN (n_0_147_1), .A (sps__n91));
NAND4_X1 i_0_147_2 (.ZN (n_0_147_0), .A1 (n_0_147_4), .A2 (n_0_147_3), .A3 (n_0_147_2), .A4 (n_0_147_1));
NAND3_X1 i_0_132_36 (.ZN (n_0_168), .A1 (n_0_132_33), .A2 (n_0_132_34), .A3 (n_0_132_35));
NAND2_X1 i_0_132_35 (.ZN (n_0_132_35), .A1 (n_0_132_24), .A2 (\mem[4][3] ));
NAND2_X1 i_0_132_34 (.ZN (n_0_132_34), .A1 (n_0_132_23), .A2 (\mem[4][3] ));
NAND3_X1 i_0_132_33 (.ZN (n_0_132_33), .A1 (n_0_132_26), .A2 (n_0_132_32), .A3 (n_0_132_29));
NOR2_X1 i_0_132_32 (.ZN (n_0_132_32), .A1 (n_0_132_0), .A2 (n_0_132_18));
INV_X1 i_0_132_31 (.ZN (n_0_132_31), .A (n_0_132_18));
INV_X1 i_0_132_30 (.ZN (n_0_132_30), .A (n_0_132_0));
NOR2_X1 i_0_132_29 (.ZN (n_0_132_29), .A1 (n_0_132_5), .A2 (n_0_132_14));
INV_X1 i_0_132_28 (.ZN (n_0_132_28), .A (n_0_132_14));
INV_X1 i_0_132_27 (.ZN (n_0_132_27), .A (n_0_132_5));
INV_X1 i_0_132_26 (.ZN (n_0_132_26), .A (n_0_132_25));
NAND2_X1 i_0_132_25 (.ZN (n_0_132_25), .A1 (n_0_132_10), .A2 (data[3]));
NAND2_X1 i_0_132_24 (.ZN (n_0_132_24), .A1 (n_0_132_30), .A2 (n_0_132_27));
NAND3_X1 i_0_132_23 (.ZN (n_0_132_23), .A1 (n_0_132_31), .A2 (n_0_132_28), .A3 (n_0_132_10));
INV_X1 i_0_132_22 (.ZN (n_0_132_22), .A (sps__n34));
INV_X1 i_0_132_21 (.ZN (n_0_132_21), .A (sps__n9));
INV_X1 i_0_132_20 (.ZN (n_0_132_20), .A (sps__n15));
INV_X1 i_0_132_19 (.ZN (n_0_132_19), .A (sps__n51));
NAND4_X1 i_0_132_18 (.ZN (n_0_132_18), .A1 (n_0_132_22), .A2 (n_0_132_21), .A3 (n_0_132_20), .A4 (n_0_132_19));
INV_X1 i_0_132_17 (.ZN (n_0_132_17), .A (sps__n63));
INV_X1 i_0_132_12 (.ZN (n_0_132_16), .A (sps__n74));
INV_X1 i_0_132_11 (.ZN (n_0_132_15), .A (sps__n86));
NAND4_X1 i_0_132_6 (.ZN (n_0_132_14), .A1 (n_0_132_17), .A2 (n_0_132_16), .A3 (n_0_132_15), .A4 (sps__n3));
INV_X1 i_0_132_5 (.ZN (n_0_132_13), .A (sps__n112));
INV_X1 i_0_132_4 (.ZN (n_0_132_12), .A (sps__n99));
NAND3_X1 i_0_132_1 (.ZN (n_0_132_11), .A1 (n_0_132_13), .A2 (n_0_132_12), .A3 (sps__n122));
INV_X1 i_0_132_0 (.ZN (n_0_132_10), .A (n_0_132_11));
INV_X1 i_0_132_16 (.ZN (n_0_132_9), .A (sps__n67));
INV_X1 i_0_132_15 (.ZN (n_0_132_8), .A (sps__n19));
INV_X1 i_0_132_14 (.ZN (n_0_132_7), .A (sps__n81));
INV_X1 i_0_132_13 (.ZN (n_0_132_6), .A (sps__n104));
NAND4_X1 i_0_132_3 (.ZN (n_0_132_5), .A1 (n_0_132_9), .A2 (n_0_132_8), .A3 (n_0_132_7), .A4 (n_0_132_6));
INV_X1 i_0_132_10 (.ZN (n_0_132_4), .A (sps__n55));
INV_X1 i_0_132_9 (.ZN (n_0_132_3), .A (sps__n28));
INV_X1 i_0_132_8 (.ZN (n_0_132_2), .A (sps__n43));
INV_X1 i_0_132_7 (.ZN (n_0_132_1), .A (sps__n92));
NAND4_X1 i_0_132_2 (.ZN (n_0_132_0), .A1 (n_0_132_4), .A2 (n_0_132_3), .A3 (n_0_132_2), .A4 (n_0_132_1));
NAND3_X1 i_0_131_36 (.ZN (n_0_167), .A1 (n_0_131_33), .A2 (n_0_131_34), .A3 (n_0_131_35));
NAND2_X1 i_0_131_35 (.ZN (n_0_131_35), .A1 (n_0_131_24), .A2 (\mem[4][4] ));
NAND2_X1 i_0_131_34 (.ZN (n_0_131_34), .A1 (n_0_131_23), .A2 (\mem[4][4] ));
NAND3_X1 i_0_131_33 (.ZN (n_0_131_33), .A1 (n_0_131_26), .A2 (n_0_131_32), .A3 (n_0_131_29));
NOR2_X1 i_0_131_32 (.ZN (n_0_131_32), .A1 (n_0_131_0), .A2 (n_0_131_18));
INV_X1 i_0_131_31 (.ZN (n_0_131_31), .A (n_0_131_18));
INV_X1 i_0_131_30 (.ZN (n_0_131_30), .A (n_0_131_0));
NOR2_X1 i_0_131_29 (.ZN (n_0_131_29), .A1 (n_0_131_5), .A2 (n_0_131_14));
INV_X1 i_0_131_28 (.ZN (n_0_131_28), .A (n_0_131_14));
INV_X1 i_0_131_27 (.ZN (n_0_131_27), .A (n_0_131_5));
INV_X1 i_0_131_26 (.ZN (n_0_131_26), .A (n_0_131_25));
NAND2_X1 i_0_131_25 (.ZN (n_0_131_25), .A1 (n_0_131_10), .A2 (data[4]));
NAND2_X1 i_0_131_24 (.ZN (n_0_131_24), .A1 (n_0_131_30), .A2 (n_0_131_27));
NAND3_X1 i_0_131_23 (.ZN (n_0_131_23), .A1 (n_0_131_31), .A2 (n_0_131_28), .A3 (n_0_131_10));
INV_X1 i_0_131_22 (.ZN (n_0_131_22), .A (sps__n34));
INV_X1 i_0_131_21 (.ZN (n_0_131_21), .A (sps__n9));
INV_X1 i_0_131_20 (.ZN (n_0_131_20), .A (sps__n15));
INV_X1 i_0_131_19 (.ZN (n_0_131_19), .A (sps__n51));
NAND4_X1 i_0_131_18 (.ZN (n_0_131_18), .A1 (n_0_131_22), .A2 (n_0_131_21), .A3 (n_0_131_20), .A4 (n_0_131_19));
INV_X1 i_0_131_17 (.ZN (n_0_131_17), .A (sps__n62));
INV_X1 i_0_131_12 (.ZN (n_0_131_16), .A (sps__n75));
INV_X1 i_0_131_11 (.ZN (n_0_131_15), .A (sps__n86));
NAND4_X1 i_0_131_6 (.ZN (n_0_131_14), .A1 (n_0_131_17), .A2 (n_0_131_16), .A3 (n_0_131_15), .A4 (sps__n3));
INV_X1 i_0_131_5 (.ZN (n_0_131_13), .A (sps__n112));
INV_X1 i_0_131_4 (.ZN (n_0_131_12), .A (sps__n99));
NAND3_X1 i_0_131_1 (.ZN (n_0_131_11), .A1 (n_0_131_13), .A2 (n_0_131_12), .A3 (sps__n122));
INV_X1 i_0_131_0 (.ZN (n_0_131_10), .A (n_0_131_11));
INV_X1 i_0_131_16 (.ZN (n_0_131_9), .A (sps__n67));
INV_X1 i_0_131_15 (.ZN (n_0_131_8), .A (sps__n19));
INV_X1 i_0_131_14 (.ZN (n_0_131_7), .A (sps__n81));
INV_X1 i_0_131_13 (.ZN (n_0_131_6), .A (sps__n105));
NAND4_X1 i_0_131_3 (.ZN (n_0_131_5), .A1 (n_0_131_9), .A2 (n_0_131_8), .A3 (n_0_131_7), .A4 (n_0_131_6));
INV_X1 i_0_131_10 (.ZN (n_0_131_4), .A (sps__n55));
INV_X1 i_0_131_9 (.ZN (n_0_131_3), .A (sps__n28));
INV_X1 i_0_131_8 (.ZN (n_0_131_2), .A (sps__n43));
INV_X1 i_0_131_7 (.ZN (n_0_131_1), .A (sps__n92));
NAND4_X1 i_0_131_2 (.ZN (n_0_131_0), .A1 (n_0_131_4), .A2 (n_0_131_3), .A3 (n_0_131_2), .A4 (n_0_131_1));
NAND3_X1 i_0_130_31 (.ZN (n_0_130_30), .A1 (n_0_130_27), .A2 (n_0_130_28), .A3 (n_0_130_29));
NOR2_X1 i_0_130_30 (.ZN (n_0_130_29), .A1 (n_0_130_13), .A2 (n_0_130_23));
NOR2_X1 i_0_130_29 (.ZN (n_0_130_28), .A1 (n_0_130_22), .A2 (n_0_130_21));
NOR2_X1 i_0_130_28 (.ZN (n_0_130_27), .A1 (n_0_130_17), .A2 (n_0_130_20));
NOR2_X1 i_0_130_27 (.ZN (n_0_130_26), .A1 (n_0_130_17), .A2 (n_0_130_13));
NOR2_X1 i_0_130_26 (.ZN (n_0_130_25), .A1 (n_0_130_20), .A2 (n_0_130_21));
NOR2_X1 i_0_130_25 (.ZN (n_0_130_24), .A1 (n_0_130_22), .A2 (n_0_130_23));
NAND3_X1 i_0_130_24 (.ZN (n_0_130_23), .A1 (n_0_130_4), .A2 (n_0_130_2), .A3 (n_0_130_6));
NAND3_X1 i_0_130_23 (.ZN (n_0_130_22), .A1 (n_0_130_1), .A2 (n_0_130_3), .A3 (n_0_130_5));
NAND3_X1 i_0_130_22 (.ZN (n_0_130_21), .A1 (n_0_130_10), .A2 (n_0_130_8), .A3 (n_0_130_12));
NAND3_X1 i_0_130_21 (.ZN (n_0_130_20), .A1 (n_0_130_7), .A2 (n_0_130_9), .A3 (n_0_130_11));
NAND2_X1 i_0_130_20 (.ZN (n_0_130_19), .A1 (n_0_130_30), .A2 (\mem[5][4] ));
INV_X1 i_0_130_19 (.ZN (n_0_130_18), .A (sps__n112));
NAND4_X1 i_0_130_18 (.ZN (n_0_130_17), .A1 (n_0_130_18), .A2 (sps__n3), .A3 (sps__n121), .A4 (sps__n99));
INV_X1 i_0_130_17 (.ZN (n_0_130_16), .A (sps__n21));
INV_X1 i_0_130_16 (.ZN (n_0_130_15), .A (sps__n80));
INV_X1 i_0_130_15 (.ZN (n_0_130_14), .A (sps__n103));
NAND3_X1 i_0_130_14 (.ZN (n_0_130_13), .A1 (n_0_130_16), .A2 (n_0_130_15), .A3 (n_0_130_14));
INV_X1 i_0_130_13 (.ZN (n_0_130_12), .A (sps__n63));
INV_X1 i_0_130_12 (.ZN (n_0_130_11), .A (sps__n74));
INV_X1 i_0_130_11 (.ZN (n_0_130_10), .A (sps__n8));
INV_X1 i_0_130_10 (.ZN (n_0_130_9), .A (sps__n14));
INV_X1 i_0_130_9 (.ZN (n_0_130_8), .A (sps__n87));
INV_X1 i_0_130_8 (.ZN (n_0_130_7), .A (sps__n35));
INV_X1 i_0_130_7 (.ZN (n_0_130_6), .A (sps__n91));
INV_X1 i_0_130_6 (.ZN (n_0_130_5), .A (sps__n67));
INV_X1 i_0_130_5 (.ZN (n_0_130_4), .A (sps__n26));
INV_X1 i_0_130_4 (.ZN (n_0_130_3), .A (sps__n44));
INV_X1 i_0_130_3 (.ZN (n_0_130_2), .A (sps__n49));
INV_X1 i_0_130_2 (.ZN (n_0_130_1), .A (sps__n57));
NAND4_X1 i_0_130_1 (.ZN (n_0_130_0), .A1 (n_0_130_26), .A2 (n_0_130_25), .A3 (n_0_130_24), .A4 (data[4]));
NAND2_X1 i_0_130_0 (.ZN (n_0_166), .A1 (n_0_130_19), .A2 (n_0_130_0));
NAND3_X1 i_0_113_31 (.ZN (n_0_113_30), .A1 (n_0_113_27), .A2 (n_0_113_28), .A3 (n_0_113_29));
NOR2_X1 i_0_113_30 (.ZN (n_0_113_29), .A1 (n_0_113_13), .A2 (n_0_113_23));
NOR2_X1 i_0_113_29 (.ZN (n_0_113_28), .A1 (n_0_113_22), .A2 (n_0_113_21));
NOR2_X1 i_0_113_28 (.ZN (n_0_113_27), .A1 (n_0_113_17), .A2 (n_0_113_20));
NOR2_X1 i_0_113_27 (.ZN (n_0_113_26), .A1 (n_0_113_17), .A2 (n_0_113_13));
NOR2_X1 i_0_113_26 (.ZN (n_0_113_25), .A1 (n_0_113_20), .A2 (n_0_113_21));
NOR2_X1 i_0_113_25 (.ZN (n_0_113_24), .A1 (n_0_113_22), .A2 (n_0_113_23));
NAND3_X1 i_0_113_24 (.ZN (n_0_113_23), .A1 (n_0_113_4), .A2 (n_0_113_2), .A3 (n_0_113_6));
NAND3_X1 i_0_113_23 (.ZN (n_0_113_22), .A1 (n_0_113_1), .A2 (n_0_113_3), .A3 (n_0_113_5));
NAND3_X1 i_0_113_22 (.ZN (n_0_113_21), .A1 (n_0_113_10), .A2 (n_0_113_8), .A3 (n_0_113_12));
NAND3_X1 i_0_113_21 (.ZN (n_0_113_20), .A1 (n_0_113_7), .A2 (n_0_113_9), .A3 (n_0_113_11));
NAND2_X1 i_0_113_20 (.ZN (n_0_113_19), .A1 (n_0_113_30), .A2 (\mem[6][4] ));
INV_X1 i_0_113_19 (.ZN (n_0_113_18), .A (sps__n99));
NAND4_X1 i_0_113_18 (.ZN (n_0_113_17), .A1 (n_0_113_18), .A2 (sps__n3), .A3 (sps__n122), .A4 (sps__n112));
INV_X1 i_0_113_17 (.ZN (n_0_113_16), .A (sps__n19));
INV_X1 i_0_113_16 (.ZN (n_0_113_15), .A (sps__n81));
INV_X1 i_0_113_15 (.ZN (n_0_113_14), .A (sps__n104));
NAND3_X1 i_0_113_14 (.ZN (n_0_113_13), .A1 (n_0_113_16), .A2 (n_0_113_15), .A3 (n_0_113_14));
INV_X1 i_0_113_13 (.ZN (n_0_113_12), .A (sps__n63));
INV_X1 i_0_113_12 (.ZN (n_0_113_11), .A (sps__n75));
INV_X1 i_0_113_11 (.ZN (n_0_113_10), .A (sps__n8));
INV_X1 i_0_113_10 (.ZN (n_0_113_9), .A (sps__n15));
INV_X1 i_0_113_9 (.ZN (n_0_113_8), .A (sps__n87));
INV_X1 i_0_113_8 (.ZN (n_0_113_7), .A (sps__n34));
INV_X1 i_0_113_7 (.ZN (n_0_113_6), .A (sps__n91));
INV_X1 i_0_113_6 (.ZN (n_0_113_5), .A (sps__n67));
INV_X1 i_0_113_5 (.ZN (n_0_113_4), .A (sps__n26));
INV_X1 i_0_113_4 (.ZN (n_0_113_3), .A (sps__n43));
INV_X1 i_0_113_3 (.ZN (n_0_113_2), .A (sps__n50));
INV_X1 i_0_113_2 (.ZN (n_0_113_1), .A (sps__n57));
NAND4_X1 i_0_113_1 (.ZN (n_0_113_0), .A1 (n_0_113_26), .A2 (n_0_113_25), .A3 (n_0_113_24), .A4 (data[4]));
NAND2_X1 i_0_113_0 (.ZN (n_0_165), .A1 (n_0_113_19), .A2 (n_0_113_0));
NAND3_X1 i_0_96_27 (.ZN (n_0_96_26), .A1 (n_0_96_23), .A2 (n_0_96_24), .A3 (n_0_96_25));
NOR2_X1 i_0_96_26 (.ZN (n_0_96_25), .A1 (n_0_96_17), .A2 (n_0_96_13));
NOR2_X1 i_0_96_25 (.ZN (n_0_96_24), .A1 (n_0_96_19), .A2 (n_0_96_20));
NOR2_X1 i_0_96_24 (.ZN (n_0_96_23), .A1 (n_0_96_21), .A2 (n_0_96_22));
NAND3_X1 i_0_96_23 (.ZN (n_0_96_22), .A1 (n_0_96_4), .A2 (n_0_96_2), .A3 (n_0_96_6));
NAND3_X1 i_0_96_22 (.ZN (n_0_96_21), .A1 (n_0_96_1), .A2 (n_0_96_3), .A3 (n_0_96_5));
NAND3_X1 i_0_96_21 (.ZN (n_0_96_20), .A1 (n_0_96_10), .A2 (n_0_96_8), .A3 (n_0_96_12));
NAND3_X1 i_0_96_20 (.ZN (n_0_96_19), .A1 (n_0_96_7), .A2 (n_0_96_9), .A3 (n_0_96_11));
NAND2_X1 i_0_96_19 (.ZN (n_0_96_18), .A1 (n_0_96_26), .A2 (\mem[7][2] ));
NAND4_X1 i_0_96_18 (.ZN (n_0_96_17), .A1 (sps__n1), .A2 (sps__n121), .A3 (sps__n112), .A4 (sps__n97));
INV_X1 i_0_96_17 (.ZN (n_0_96_16), .A (sps__n21));
INV_X1 i_0_96_16 (.ZN (n_0_96_15), .A (sps__n80));
INV_X1 i_0_96_15 (.ZN (n_0_96_14), .A (sps__n103));
NAND3_X1 i_0_96_14 (.ZN (n_0_96_13), .A1 (n_0_96_16), .A2 (n_0_96_15), .A3 (n_0_96_14));
INV_X1 i_0_96_13 (.ZN (n_0_96_12), .A (sps__n63));
INV_X1 i_0_96_12 (.ZN (n_0_96_11), .A (sps__n75));
INV_X1 i_0_96_11 (.ZN (n_0_96_10), .A (sps__n8));
INV_X1 i_0_96_10 (.ZN (n_0_96_9), .A (sps__n13));
INV_X1 i_0_96_9 (.ZN (n_0_96_8), .A (sps__n87));
INV_X1 i_0_96_8 (.ZN (n_0_96_7), .A (sps__n35));
INV_X1 i_0_96_7 (.ZN (n_0_96_6), .A (sps__n93));
INV_X1 i_0_96_6 (.ZN (n_0_96_5), .A (sps__n67));
INV_X1 i_0_96_5 (.ZN (n_0_96_4), .A (sps__n27));
INV_X1 i_0_96_4 (.ZN (n_0_96_3), .A (sps__n44));
INV_X1 i_0_96_3 (.ZN (n_0_96_2), .A (sps__n49));
INV_X1 i_0_96_2 (.ZN (n_0_96_1), .A (sps__n57));
NAND4_X1 i_0_96_1 (.ZN (n_0_96_0), .A1 (n_0_96_25), .A2 (n_0_96_24), .A3 (n_0_96_23), .A4 (data[2]));
NAND2_X1 i_0_96_0 (.ZN (n_0_164), .A1 (n_0_96_18), .A2 (n_0_96_0));
NAND3_X1 i_0_81_27 (.ZN (n_0_81_26), .A1 (n_0_81_23), .A2 (n_0_81_24), .A3 (n_0_81_25));
NOR2_X1 i_0_81_26 (.ZN (n_0_81_25), .A1 (n_0_81_17), .A2 (n_0_81_13));
NOR2_X1 i_0_81_25 (.ZN (n_0_81_24), .A1 (n_0_81_19), .A2 (n_0_81_20));
NOR2_X1 i_0_81_24 (.ZN (n_0_81_23), .A1 (n_0_81_21), .A2 (n_0_81_22));
NAND3_X1 i_0_81_23 (.ZN (n_0_81_22), .A1 (n_0_81_4), .A2 (n_0_81_2), .A3 (n_0_81_6));
NAND3_X1 i_0_81_22 (.ZN (n_0_81_21), .A1 (n_0_81_1), .A2 (n_0_81_3), .A3 (n_0_81_5));
NAND3_X1 i_0_81_21 (.ZN (n_0_81_20), .A1 (n_0_81_10), .A2 (n_0_81_8), .A3 (n_0_81_12));
NAND3_X1 i_0_81_20 (.ZN (n_0_81_19), .A1 (n_0_81_7), .A2 (n_0_81_9), .A3 (n_0_81_11));
NAND2_X1 i_0_81_19 (.ZN (n_0_81_18), .A1 (n_0_81_26), .A2 (\mem[7][3] ));
NAND4_X1 i_0_81_18 (.ZN (n_0_81_17), .A1 (sps__n1), .A2 (sps__n121), .A3 (sps__n114), .A4 (sps__n97));
INV_X1 i_0_81_17 (.ZN (n_0_81_16), .A (sps__n21));
INV_X1 i_0_81_16 (.ZN (n_0_81_15), .A (sps__n80));
INV_X1 i_0_81_15 (.ZN (n_0_81_14), .A (sps__n103));
NAND3_X1 i_0_81_14 (.ZN (n_0_81_13), .A1 (n_0_81_16), .A2 (n_0_81_15), .A3 (n_0_81_14));
INV_X1 i_0_81_13 (.ZN (n_0_81_12), .A (sps__n61));
INV_X1 i_0_81_12 (.ZN (n_0_81_11), .A (sps__n74));
INV_X1 i_0_81_11 (.ZN (n_0_81_10), .A (sps__n8));
INV_X1 i_0_81_10 (.ZN (n_0_81_9), .A (sps__n13));
INV_X1 i_0_81_9 (.ZN (n_0_81_8), .A (sps__n85));
INV_X1 i_0_81_8 (.ZN (n_0_81_7), .A (sps__n36));
INV_X1 i_0_81_7 (.ZN (n_0_81_6), .A (sps__n91));
INV_X1 i_0_81_6 (.ZN (n_0_81_5), .A (sps__n68));
INV_X1 i_0_81_5 (.ZN (n_0_81_4), .A (sps__n26));
INV_X1 i_0_81_4 (.ZN (n_0_81_3), .A (sps__n44));
INV_X1 i_0_81_3 (.ZN (n_0_81_2), .A (sps__n49));
INV_X1 i_0_81_2 (.ZN (n_0_81_1), .A (sps__n55));
NAND4_X1 i_0_81_1 (.ZN (n_0_81_0), .A1 (n_0_81_25), .A2 (n_0_81_24), .A3 (n_0_81_23), .A4 (data[3]));
NAND2_X1 i_0_81_0 (.ZN (n_0_163), .A1 (n_0_81_18), .A2 (n_0_81_0));
NAND3_X1 i_0_80_27 (.ZN (n_0_80_26), .A1 (n_0_80_23), .A2 (n_0_80_24), .A3 (n_0_80_25));
NOR2_X1 i_0_80_26 (.ZN (n_0_80_25), .A1 (n_0_80_17), .A2 (n_0_80_13));
NOR2_X1 i_0_80_25 (.ZN (n_0_80_24), .A1 (n_0_80_19), .A2 (n_0_80_20));
NOR2_X1 i_0_80_24 (.ZN (n_0_80_23), .A1 (n_0_80_21), .A2 (n_0_80_22));
NAND3_X1 i_0_80_23 (.ZN (n_0_80_22), .A1 (n_0_80_4), .A2 (n_0_80_2), .A3 (n_0_80_6));
NAND3_X1 i_0_80_22 (.ZN (n_0_80_21), .A1 (n_0_80_1), .A2 (n_0_80_3), .A3 (n_0_80_5));
NAND3_X1 i_0_80_21 (.ZN (n_0_80_20), .A1 (n_0_80_10), .A2 (n_0_80_8), .A3 (n_0_80_12));
NAND3_X1 i_0_80_20 (.ZN (n_0_80_19), .A1 (n_0_80_7), .A2 (n_0_80_9), .A3 (n_0_80_11));
NAND2_X1 i_0_80_19 (.ZN (n_0_80_18), .A1 (n_0_80_26), .A2 (\mem[7][4] ));
NAND4_X1 i_0_80_18 (.ZN (n_0_80_17), .A1 (sps__n3), .A2 (sps__n121), .A3 (sps__n114), .A4 (sps__n97));
INV_X1 i_0_80_17 (.ZN (n_0_80_16), .A (sps__n21));
INV_X1 i_0_80_16 (.ZN (n_0_80_15), .A (sps__n80));
INV_X1 i_0_80_15 (.ZN (n_0_80_14), .A (sps__n103));
NAND3_X1 i_0_80_14 (.ZN (n_0_80_13), .A1 (n_0_80_16), .A2 (n_0_80_15), .A3 (n_0_80_14));
INV_X1 i_0_80_13 (.ZN (n_0_80_12), .A (sps__n61));
INV_X1 i_0_80_12 (.ZN (n_0_80_11), .A (sps__n74));
INV_X1 i_0_80_11 (.ZN (n_0_80_10), .A (sps__n8));
INV_X1 i_0_80_10 (.ZN (n_0_80_9), .A (sps__n13));
INV_X1 i_0_80_9 (.ZN (n_0_80_8), .A (sps__n87));
INV_X1 i_0_80_8 (.ZN (n_0_80_7), .A (sps__n36));
INV_X1 i_0_80_7 (.ZN (n_0_80_6), .A (sps__n91));
INV_X1 i_0_80_6 (.ZN (n_0_80_5), .A (sps__n68));
INV_X1 i_0_80_5 (.ZN (n_0_80_4), .A (sps__n26));
INV_X1 i_0_80_4 (.ZN (n_0_80_3), .A (sps__n44));
INV_X1 i_0_80_3 (.ZN (n_0_80_2), .A (sps__n49));
INV_X1 i_0_80_2 (.ZN (n_0_80_1), .A (sps__n55));
NAND4_X1 i_0_80_1 (.ZN (n_0_80_0), .A1 (n_0_80_25), .A2 (n_0_80_24), .A3 (n_0_80_23), .A4 (data[4]));
NAND2_X1 i_0_80_0 (.ZN (n_0_162), .A1 (n_0_80_18), .A2 (n_0_80_0));
NAND3_X1 i_0_79_35 (.ZN (n_0_161), .A1 (n_0_79_32), .A2 (n_0_79_33), .A3 (n_0_79_34));
NAND2_X1 i_0_79_34 (.ZN (n_0_79_34), .A1 (n_0_79_23), .A2 (\mem[8][3] ));
NAND3_X1 i_0_79_29 (.ZN (n_0_79_33), .A1 (n_0_79_26), .A2 (n_0_79_31), .A3 (n_0_79_28));
NAND2_X1 i_0_79_28 (.ZN (n_0_79_32), .A1 (n_0_79_27), .A2 (\mem[8][3] ));
NOR2_X1 i_0_79_24 (.ZN (n_0_79_31), .A1 (n_0_79_18), .A2 (n_0_79_0));
INV_X1 i_0_79_23 (.ZN (n_0_79_30), .A (n_0_79_0));
INV_X1 i_0_79_22 (.ZN (n_0_79_29), .A (n_0_79_18));
INV_X1 i_0_79_21 (.ZN (n_0_79_28), .A (n_0_79_5));
NAND3_X1 i_0_79_20 (.ZN (n_0_79_27), .A1 (n_0_79_28), .A2 (n_0_79_30), .A3 (n_0_79_9));
NOR2_X1 i_0_79_19 (.ZN (n_0_79_26), .A1 (n_0_79_14), .A2 (n_0_79_24));
INV_X1 i_0_79_18 (.ZN (n_0_79_25), .A (n_0_79_14));
NAND2_X1 i_0_79_17 (.ZN (n_0_79_24), .A1 (n_0_79_9), .A2 (data[3]));
NAND2_X1 i_0_79_16 (.ZN (n_0_79_23), .A1 (n_0_79_29), .A2 (n_0_79_25));
INV_X1 i_0_79_33 (.ZN (n_0_79_22), .A (sps__n34));
INV_X1 i_0_79_32 (.ZN (n_0_79_21), .A (sps__n8));
INV_X1 i_0_79_31 (.ZN (n_0_79_20), .A (sps__n14));
INV_X1 i_0_79_30 (.ZN (n_0_79_19), .A (sps__n50));
NAND4_X1 i_0_79_3 (.ZN (n_0_79_18), .A1 (n_0_79_22), .A2 (n_0_79_21), .A3 (n_0_79_20), .A4 (n_0_79_19));
INV_X1 i_0_79_27 (.ZN (n_0_79_17), .A (sps__n62));
INV_X1 i_0_79_26 (.ZN (n_0_79_16), .A (sps__n74));
INV_X1 i_0_79_25 (.ZN (n_0_79_15), .A (sps__n85));
NAND4_X1 i_0_79_8 (.ZN (n_0_79_14), .A1 (n_0_79_17), .A2 (n_0_79_16), .A3 (n_0_79_15), .A4 (sps__n3));
INV_X1 i_0_79_15 (.ZN (n_0_79_13), .A (sps__n121));
INV_X1 i_0_79_14 (.ZN (n_0_79_12), .A (sps__n112));
INV_X1 i_0_79_13 (.ZN (n_0_79_11), .A (sps__n99));
NAND3_X1 i_0_79_12 (.ZN (n_0_79_10), .A1 (n_0_79_13), .A2 (n_0_79_12), .A3 (n_0_79_11));
INV_X1 i_0_79_11 (.ZN (n_0_79_9), .A (n_0_79_10));
INV_X1 i_0_79_10 (.ZN (n_0_79_8), .A (sps__n68));
INV_X1 i_0_79_9 (.ZN (n_0_79_7), .A (sps__n19));
INV_X1 i_0_79_7 (.ZN (n_0_79_6), .A (sps__n81));
NAND4_X1 i_0_79_6 (.ZN (n_0_79_5), .A1 (n_0_79_8), .A2 (n_0_79_7), .A3 (n_0_79_6), .A4 (sps__n104));
INV_X1 i_0_79_5 (.ZN (n_0_79_4), .A (sps__n55));
INV_X1 i_0_79_4 (.ZN (n_0_79_3), .A (sps__n28));
INV_X1 i_0_79_2 (.ZN (n_0_79_2), .A (sps__n44));
INV_X1 i_0_79_1 (.ZN (n_0_79_1), .A (sps__n91));
NAND4_X1 i_0_79_0 (.ZN (n_0_79_0), .A1 (n_0_79_4), .A2 (n_0_79_3), .A3 (n_0_79_2), .A4 (n_0_79_1));
NAND3_X1 i_0_63_35 (.ZN (n_0_160), .A1 (n_0_63_32), .A2 (n_0_63_33), .A3 (n_0_63_34));
NAND2_X1 i_0_63_34 (.ZN (n_0_63_34), .A1 (n_0_63_23), .A2 (\mem[8][4] ));
NAND3_X1 i_0_63_29 (.ZN (n_0_63_33), .A1 (n_0_63_26), .A2 (n_0_63_31), .A3 (n_0_63_28));
NAND2_X1 i_0_63_28 (.ZN (n_0_63_32), .A1 (n_0_63_27), .A2 (\mem[8][4] ));
NOR2_X1 i_0_63_24 (.ZN (n_0_63_31), .A1 (n_0_63_18), .A2 (n_0_63_0));
INV_X1 i_0_63_23 (.ZN (n_0_63_30), .A (n_0_63_0));
INV_X1 i_0_63_22 (.ZN (n_0_63_29), .A (n_0_63_18));
INV_X1 i_0_63_21 (.ZN (n_0_63_28), .A (n_0_63_5));
NAND3_X1 i_0_63_20 (.ZN (n_0_63_27), .A1 (n_0_63_28), .A2 (n_0_63_30), .A3 (n_0_63_9));
NOR2_X1 i_0_63_19 (.ZN (n_0_63_26), .A1 (n_0_63_14), .A2 (n_0_63_24));
INV_X1 i_0_63_18 (.ZN (n_0_63_25), .A (n_0_63_14));
NAND2_X1 i_0_63_17 (.ZN (n_0_63_24), .A1 (n_0_63_9), .A2 (data[4]));
NAND2_X1 i_0_63_16 (.ZN (n_0_63_23), .A1 (n_0_63_29), .A2 (n_0_63_25));
INV_X1 i_0_63_33 (.ZN (n_0_63_22), .A (sps__n34));
INV_X1 i_0_63_32 (.ZN (n_0_63_21), .A (sps__n8));
INV_X1 i_0_63_31 (.ZN (n_0_63_20), .A (sps__n14));
INV_X1 i_0_63_30 (.ZN (n_0_63_19), .A (sps__n50));
NAND4_X1 i_0_63_3 (.ZN (n_0_63_18), .A1 (n_0_63_22), .A2 (n_0_63_21), .A3 (n_0_63_20), .A4 (n_0_63_19));
INV_X1 i_0_63_27 (.ZN (n_0_63_17), .A (sps__n63));
INV_X1 i_0_63_26 (.ZN (n_0_63_16), .A (sps__n74));
INV_X1 i_0_63_25 (.ZN (n_0_63_15), .A (sps__n87));
NAND4_X1 i_0_63_8 (.ZN (n_0_63_14), .A1 (n_0_63_17), .A2 (n_0_63_16), .A3 (n_0_63_15), .A4 (sps__n3));
INV_X1 i_0_63_15 (.ZN (n_0_63_13), .A (sps__n122));
INV_X1 i_0_63_14 (.ZN (n_0_63_12), .A (sps__n112));
INV_X1 i_0_63_13 (.ZN (n_0_63_11), .A (sps__n99));
NAND3_X1 i_0_63_12 (.ZN (n_0_63_10), .A1 (n_0_63_13), .A2 (n_0_63_12), .A3 (n_0_63_11));
INV_X1 i_0_63_11 (.ZN (n_0_63_9), .A (n_0_63_10));
INV_X1 i_0_63_10 (.ZN (n_0_63_8), .A (sps__n67));
INV_X1 i_0_63_9 (.ZN (n_0_63_7), .A (sps__n19));
INV_X1 i_0_63_7 (.ZN (n_0_63_6), .A (sps__n81));
NAND4_X1 i_0_63_6 (.ZN (n_0_63_5), .A1 (n_0_63_8), .A2 (n_0_63_7), .A3 (n_0_63_6), .A4 (sps__n104));
INV_X1 i_0_63_5 (.ZN (n_0_63_4), .A (sps__n57));
INV_X1 i_0_63_4 (.ZN (n_0_63_3), .A (sps__n26));
INV_X1 i_0_63_2 (.ZN (n_0_63_2), .A (sps__n43));
INV_X1 i_0_63_1 (.ZN (n_0_63_1), .A (sps__n91));
NAND4_X1 i_0_63_0 (.ZN (n_0_63_0), .A1 (n_0_63_4), .A2 (n_0_63_3), .A3 (n_0_63_2), .A4 (n_0_63_1));
NOR2_X1 i_0_62_34 (.ZN (n_0_62_33), .A1 (n_0_62_19), .A2 (n_0_62_0));
INV_X1 i_0_62_33 (.ZN (n_0_62_32), .A (n_0_62_0));
INV_X1 i_0_62_28 (.ZN (n_0_62_31), .A (n_0_62_19));
NAND2_X1 i_0_62_27 (.ZN (n_0_62_30), .A1 (n_0_62_29), .A2 (\mem[9][4] ));
NAND3_X1 i_0_62_23 (.ZN (n_0_62_29), .A1 (n_0_62_5), .A2 (n_0_62_32), .A3 (n_0_62_10));
NAND3_X1 i_0_62_22 (.ZN (n_0_62_28), .A1 (n_0_62_27), .A2 (n_0_62_33), .A3 (n_0_62_14));
NOR2_X1 i_0_62_21 (.ZN (n_0_62_27), .A1 (n_0_62_6), .A2 (n_0_62_26));
NAND2_X1 i_0_62_20 (.ZN (n_0_62_26), .A1 (n_0_62_10), .A2 (data[4]));
NAND2_X1 i_0_62_19 (.ZN (n_0_62_25), .A1 (n_0_62_31), .A2 (n_0_62_14));
NAND3_X1 i_0_62_18 (.ZN (n_0_159), .A1 (n_0_62_28), .A2 (n_0_62_30), .A3 (n_0_62_24));
NAND2_X1 i_0_62_17 (.ZN (n_0_62_24), .A1 (n_0_62_25), .A2 (\mem[9][4] ));
INV_X1 i_0_62_32 (.ZN (n_0_62_23), .A (sps__n34));
INV_X1 i_0_62_31 (.ZN (n_0_62_22), .A (sps__n8));
INV_X1 i_0_62_30 (.ZN (n_0_62_21), .A (sps__n14));
INV_X1 i_0_62_29 (.ZN (n_0_62_20), .A (sps__n50));
NAND4_X1 i_0_62_3 (.ZN (n_0_62_19), .A1 (n_0_62_23), .A2 (n_0_62_22), .A3 (n_0_62_21), .A4 (n_0_62_20));
INV_X1 i_0_62_26 (.ZN (n_0_62_18), .A (sps__n63));
INV_X1 i_0_62_25 (.ZN (n_0_62_17), .A (sps__n74));
INV_X1 i_0_62_24 (.ZN (n_0_62_16), .A (sps__n87));
NAND4_X1 i_0_62_6 (.ZN (n_0_62_15), .A1 (n_0_62_18), .A2 (n_0_62_17), .A3 (n_0_62_16), .A4 (sps__n3));
INV_X1 i_0_62_16 (.ZN (n_0_62_14), .A (n_0_62_15));
INV_X1 i_0_62_15 (.ZN (n_0_62_13), .A (sps__n121));
INV_X1 i_0_62_14 (.ZN (n_0_62_12), .A (sps__n112));
NAND3_X1 i_0_62_13 (.ZN (n_0_62_11), .A1 (n_0_62_13), .A2 (n_0_62_12), .A3 (sps__n99));
INV_X1 i_0_62_12 (.ZN (n_0_62_10), .A (n_0_62_11));
INV_X1 i_0_62_11 (.ZN (n_0_62_9), .A (sps__n67));
INV_X1 i_0_62_10 (.ZN (n_0_62_8), .A (sps__n19));
INV_X1 i_0_62_9 (.ZN (n_0_62_7), .A (sps__n81));
NAND4_X1 i_0_62_8 (.ZN (n_0_62_6), .A1 (n_0_62_9), .A2 (n_0_62_8), .A3 (n_0_62_7), .A4 (sps__n104));
INV_X1 i_0_62_7 (.ZN (n_0_62_5), .A (n_0_62_6));
INV_X1 i_0_62_5 (.ZN (n_0_62_4), .A (sps__n57));
INV_X1 i_0_62_4 (.ZN (n_0_62_3), .A (sps__n26));
INV_X1 i_0_62_2 (.ZN (n_0_62_2), .A (sps__n43));
INV_X1 i_0_62_1 (.ZN (n_0_62_1), .A (sps__n91));
NAND4_X1 i_0_62_0 (.ZN (n_0_62_0), .A1 (n_0_62_4), .A2 (n_0_62_3), .A3 (n_0_62_2), .A4 (n_0_62_1));
NOR2_X1 i_0_45_34 (.ZN (n_0_45_33), .A1 (n_0_45_19), .A2 (n_0_45_0));
INV_X1 i_0_45_33 (.ZN (n_0_45_32), .A (n_0_45_0));
INV_X1 i_0_45_28 (.ZN (n_0_45_31), .A (n_0_45_19));
NAND2_X1 i_0_45_27 (.ZN (n_0_45_30), .A1 (n_0_45_29), .A2 (\mem[10][4] ));
NAND3_X1 i_0_45_23 (.ZN (n_0_45_29), .A1 (n_0_45_5), .A2 (n_0_45_32), .A3 (n_0_45_10));
NAND3_X1 i_0_45_22 (.ZN (n_0_45_28), .A1 (n_0_45_27), .A2 (n_0_45_33), .A3 (n_0_45_14));
NOR2_X1 i_0_45_21 (.ZN (n_0_45_27), .A1 (n_0_45_6), .A2 (n_0_45_26));
NAND2_X1 i_0_45_20 (.ZN (n_0_45_26), .A1 (n_0_45_10), .A2 (data[4]));
NAND2_X1 i_0_45_19 (.ZN (n_0_45_25), .A1 (n_0_45_31), .A2 (n_0_45_14));
NAND3_X1 i_0_45_18 (.ZN (n_0_158), .A1 (n_0_45_28), .A2 (n_0_45_30), .A3 (n_0_45_24));
NAND2_X1 i_0_45_17 (.ZN (n_0_45_24), .A1 (n_0_45_25), .A2 (\mem[10][4] ));
INV_X1 i_0_45_32 (.ZN (n_0_45_23), .A (sps__n34));
INV_X1 i_0_45_31 (.ZN (n_0_45_22), .A (sps__n8));
INV_X1 i_0_45_30 (.ZN (n_0_45_21), .A (sps__n14));
INV_X1 i_0_45_29 (.ZN (n_0_45_20), .A (sps__n50));
NAND4_X1 i_0_45_3 (.ZN (n_0_45_19), .A1 (n_0_45_23), .A2 (n_0_45_22), .A3 (n_0_45_21), .A4 (n_0_45_20));
INV_X1 i_0_45_26 (.ZN (n_0_45_18), .A (sps__n63));
INV_X1 i_0_45_25 (.ZN (n_0_45_17), .A (sps__n74));
INV_X1 i_0_45_24 (.ZN (n_0_45_16), .A (sps__n87));
NAND4_X1 i_0_45_6 (.ZN (n_0_45_15), .A1 (n_0_45_18), .A2 (n_0_45_17), .A3 (n_0_45_16), .A4 (sps__n3));
INV_X1 i_0_45_16 (.ZN (n_0_45_14), .A (n_0_45_15));
INV_X1 i_0_45_15 (.ZN (n_0_45_13), .A (sps__n122));
INV_X1 i_0_45_14 (.ZN (n_0_45_12), .A (sps__n99));
NAND3_X1 i_0_45_13 (.ZN (n_0_45_11), .A1 (n_0_45_13), .A2 (n_0_45_12), .A3 (sps__n112));
INV_X1 i_0_45_12 (.ZN (n_0_45_10), .A (n_0_45_11));
INV_X1 i_0_45_11 (.ZN (n_0_45_9), .A (sps__n67));
INV_X1 i_0_45_10 (.ZN (n_0_45_8), .A (sps__n19));
INV_X1 i_0_45_9 (.ZN (n_0_45_7), .A (sps__n81));
NAND4_X1 i_0_45_8 (.ZN (n_0_45_6), .A1 (n_0_45_9), .A2 (n_0_45_8), .A3 (n_0_45_7), .A4 (sps__n104));
INV_X1 i_0_45_7 (.ZN (n_0_45_5), .A (n_0_45_6));
INV_X1 i_0_45_5 (.ZN (n_0_45_4), .A (sps__n57));
INV_X1 i_0_45_4 (.ZN (n_0_45_3), .A (sps__n26));
INV_X1 i_0_45_2 (.ZN (n_0_45_2), .A (sps__n43));
INV_X1 i_0_45_1 (.ZN (n_0_45_1), .A (sps__n91));
NAND4_X1 i_0_45_0 (.ZN (n_0_45_0), .A1 (n_0_45_4), .A2 (n_0_45_3), .A3 (n_0_45_2), .A4 (n_0_45_1));
NAND3_X1 i_0_28_37 (.ZN (n_0_157), .A1 (n_0_28_34), .A2 (n_0_28_35), .A3 (n_0_28_36));
NAND2_X1 i_0_28_36 (.ZN (n_0_28_36), .A1 (n_0_28_25), .A2 (\mem[0][5] ));
NAND3_X1 i_0_28_35 (.ZN (n_0_28_35), .A1 (n_0_28_27), .A2 (n_0_28_33), .A3 (n_0_28_30));
NAND2_X1 i_0_28_34 (.ZN (n_0_28_34), .A1 (n_0_28_24), .A2 (\mem[0][5] ));
NOR2_X1 i_0_28_33 (.ZN (n_0_28_33), .A1 (n_0_28_0), .A2 (n_0_28_19));
INV_X1 i_0_28_32 (.ZN (n_0_28_32), .A (n_0_28_19));
INV_X1 i_0_28_31 (.ZN (n_0_28_31), .A (n_0_28_0));
NOR2_X1 i_0_28_30 (.ZN (n_0_28_30), .A1 (n_0_28_5), .A2 (n_0_28_15));
INV_X1 i_0_28_29 (.ZN (n_0_28_29), .A (n_0_28_15));
INV_X1 i_0_28_28 (.ZN (n_0_28_28), .A (n_0_28_5));
INV_X1 i_0_28_27 (.ZN (n_0_28_27), .A (n_0_28_26));
NAND2_X1 i_0_28_26 (.ZN (n_0_28_26), .A1 (n_0_28_10), .A2 (data[5]));
NAND2_X1 i_0_28_25 (.ZN (n_0_28_25), .A1 (n_0_28_31), .A2 (n_0_28_28));
NAND3_X1 i_0_28_24 (.ZN (n_0_28_24), .A1 (n_0_28_32), .A2 (n_0_28_29), .A3 (n_0_28_10));
INV_X1 i_0_28_23 (.ZN (n_0_28_23), .A (address[14]));
INV_X1 i_0_28_22 (.ZN (n_0_28_22), .A (sps__n9));
INV_X1 i_0_28_21 (.ZN (n_0_28_21), .A (sps__n15));
INV_X1 i_0_28_20 (.ZN (n_0_28_20), .A (sps__n51));
NAND4_X1 i_0_28_19 (.ZN (n_0_28_19), .A1 (n_0_28_23), .A2 (n_0_28_22), .A3 (n_0_28_21), .A4 (n_0_28_20));
INV_X1 i_0_28_18 (.ZN (n_0_28_18), .A (sps__n62));
INV_X1 i_0_28_17 (.ZN (n_0_28_17), .A (sps__n75));
INV_X1 i_0_28_12 (.ZN (n_0_28_16), .A (sps__n86));
NAND4_X1 i_0_28_11 (.ZN (n_0_28_15), .A1 (n_0_28_18), .A2 (n_0_28_17), .A3 (n_0_28_16), .A4 (sps__n2));
INV_X1 i_0_28_6 (.ZN (n_0_28_14), .A (sps__n123));
INV_X1 i_0_28_5 (.ZN (n_0_28_13), .A (sps__n112));
INV_X1 i_0_28_4 (.ZN (n_0_28_12), .A (sps__n99));
NAND3_X1 i_0_28_1 (.ZN (n_0_28_11), .A1 (n_0_28_14), .A2 (n_0_28_13), .A3 (n_0_28_12));
INV_X1 i_0_28_0 (.ZN (n_0_28_10), .A (n_0_28_11));
INV_X1 i_0_28_16 (.ZN (n_0_28_9), .A (sps__n68));
INV_X1 i_0_28_15 (.ZN (n_0_28_8), .A (address[5]));
INV_X1 i_0_28_14 (.ZN (n_0_28_7), .A (sps__n81));
INV_X1 i_0_28_13 (.ZN (n_0_28_6), .A (sps__n105));
NAND4_X1 i_0_28_3 (.ZN (n_0_28_5), .A1 (n_0_28_9), .A2 (n_0_28_8), .A3 (n_0_28_7), .A4 (n_0_28_6));
INV_X1 i_0_28_10 (.ZN (n_0_28_4), .A (sps__n55));
INV_X1 i_0_28_9 (.ZN (n_0_28_3), .A (sps__n25));
INV_X1 i_0_28_8 (.ZN (n_0_28_2), .A (sps__n42));
INV_X1 i_0_28_7 (.ZN (n_0_28_1), .A (sps__n92));
NAND4_X1 i_0_28_2 (.ZN (n_0_28_0), .A1 (n_0_28_4), .A2 (n_0_28_3), .A3 (n_0_28_2), .A4 (n_0_28_1));
NAND3_X1 i_0_152_36 (.ZN (n_0_156), .A1 (n_0_152_33), .A2 (n_0_152_34), .A3 (n_0_152_35));
NAND2_X1 i_0_152_35 (.ZN (n_0_152_35), .A1 (n_0_152_24), .A2 (\mem[1][5] ));
NAND2_X1 i_0_152_34 (.ZN (n_0_152_34), .A1 (n_0_152_23), .A2 (\mem[1][5] ));
NAND3_X1 i_0_152_33 (.ZN (n_0_152_33), .A1 (n_0_152_26), .A2 (n_0_152_32), .A3 (n_0_152_29));
NOR2_X1 i_0_152_32 (.ZN (n_0_152_32), .A1 (n_0_152_0), .A2 (n_0_152_18));
INV_X1 i_0_152_31 (.ZN (n_0_152_31), .A (n_0_152_18));
INV_X1 i_0_152_30 (.ZN (n_0_152_30), .A (n_0_152_0));
NOR2_X1 i_0_152_29 (.ZN (n_0_152_29), .A1 (n_0_152_5), .A2 (n_0_152_14));
INV_X1 i_0_152_28 (.ZN (n_0_152_28), .A (n_0_152_14));
INV_X1 i_0_152_27 (.ZN (n_0_152_27), .A (n_0_152_5));
INV_X1 i_0_152_26 (.ZN (n_0_152_26), .A (n_0_152_25));
NAND2_X1 i_0_152_25 (.ZN (n_0_152_25), .A1 (n_0_152_10), .A2 (data[5]));
NAND2_X1 i_0_152_24 (.ZN (n_0_152_24), .A1 (n_0_152_30), .A2 (n_0_152_27));
NAND3_X1 i_0_152_23 (.ZN (n_0_152_23), .A1 (n_0_152_31), .A2 (n_0_152_28), .A3 (n_0_152_10));
INV_X1 i_0_152_22 (.ZN (n_0_152_22), .A (sps__n36));
INV_X1 i_0_152_21 (.ZN (n_0_152_21), .A (sps__n7));
INV_X1 i_0_152_20 (.ZN (n_0_152_20), .A (sps__n14));
INV_X1 i_0_152_19 (.ZN (n_0_152_19), .A (sps__n51));
NAND4_X1 i_0_152_18 (.ZN (n_0_152_18), .A1 (n_0_152_22), .A2 (n_0_152_21), .A3 (n_0_152_20), .A4 (n_0_152_19));
INV_X1 i_0_152_17 (.ZN (n_0_152_17), .A (sps__n62));
INV_X1 i_0_152_12 (.ZN (n_0_152_16), .A (sps__n74));
INV_X1 i_0_152_11 (.ZN (n_0_152_15), .A (sps__n86));
NAND4_X1 i_0_152_6 (.ZN (n_0_152_14), .A1 (n_0_152_17), .A2 (n_0_152_16), .A3 (n_0_152_15), .A4 (sps__n2));
INV_X1 i_0_152_5 (.ZN (n_0_152_13), .A (sps__n123));
INV_X1 i_0_152_4 (.ZN (n_0_152_12), .A (sps__n112));
NAND3_X1 i_0_152_1 (.ZN (n_0_152_11), .A1 (n_0_152_13), .A2 (n_0_152_12), .A3 (sps__n98));
INV_X1 i_0_152_0 (.ZN (n_0_152_10), .A (n_0_152_11));
INV_X1 i_0_152_16 (.ZN (n_0_152_9), .A (sps__n68));
INV_X1 i_0_152_15 (.ZN (n_0_152_8), .A (address[5]));
INV_X1 i_0_152_14 (.ZN (n_0_152_7), .A (address[4]));
INV_X1 i_0_152_13 (.ZN (n_0_152_6), .A (sps__n103));
NAND4_X1 i_0_152_3 (.ZN (n_0_152_5), .A1 (n_0_152_9), .A2 (n_0_152_8), .A3 (n_0_152_7), .A4 (n_0_152_6));
INV_X1 i_0_152_10 (.ZN (n_0_152_4), .A (sps__n55));
INV_X1 i_0_152_9 (.ZN (n_0_152_3), .A (sps__n25));
INV_X1 i_0_152_8 (.ZN (n_0_152_2), .A (sps__n42));
INV_X1 i_0_152_7 (.ZN (n_0_152_1), .A (sps__n92));
NAND4_X1 i_0_152_2 (.ZN (n_0_152_0), .A1 (n_0_152_4), .A2 (n_0_152_3), .A3 (n_0_152_2), .A4 (n_0_152_1));
NAND3_X1 i_0_180_36 (.ZN (n_0_155), .A1 (n_0_180_33), .A2 (n_0_180_34), .A3 (n_0_180_35));
NAND2_X1 i_0_180_35 (.ZN (n_0_180_35), .A1 (n_0_180_24), .A2 (\mem[2][5] ));
NAND2_X1 i_0_180_34 (.ZN (n_0_180_34), .A1 (n_0_180_23), .A2 (\mem[2][5] ));
NAND3_X1 i_0_180_33 (.ZN (n_0_180_33), .A1 (n_0_180_26), .A2 (n_0_180_32), .A3 (n_0_180_29));
NOR2_X1 i_0_180_32 (.ZN (n_0_180_32), .A1 (n_0_180_0), .A2 (n_0_180_18));
INV_X1 i_0_180_31 (.ZN (n_0_180_31), .A (n_0_180_18));
INV_X1 i_0_180_30 (.ZN (n_0_180_30), .A (n_0_180_0));
NOR2_X1 i_0_180_29 (.ZN (n_0_180_29), .A1 (n_0_180_5), .A2 (n_0_180_14));
INV_X1 i_0_180_28 (.ZN (n_0_180_28), .A (n_0_180_14));
INV_X1 i_0_180_27 (.ZN (n_0_180_27), .A (n_0_180_5));
INV_X1 i_0_180_26 (.ZN (n_0_180_26), .A (n_0_180_25));
NAND2_X1 i_0_180_25 (.ZN (n_0_180_25), .A1 (n_0_180_10), .A2 (data[5]));
NAND2_X1 i_0_180_24 (.ZN (n_0_180_24), .A1 (n_0_180_30), .A2 (n_0_180_27));
NAND3_X1 i_0_180_23 (.ZN (n_0_180_23), .A1 (n_0_180_31), .A2 (n_0_180_28), .A3 (n_0_180_10));
INV_X1 i_0_180_22 (.ZN (n_0_180_22), .A (sps__n36));
INV_X1 i_0_180_21 (.ZN (n_0_180_21), .A (sps__n7));
INV_X1 i_0_180_20 (.ZN (n_0_180_20), .A (sps__n15));
INV_X1 i_0_180_19 (.ZN (n_0_180_19), .A (sps__n51));
NAND4_X1 i_0_180_18 (.ZN (n_0_180_18), .A1 (n_0_180_22), .A2 (n_0_180_21), .A3 (n_0_180_20), .A4 (n_0_180_19));
INV_X1 i_0_180_17 (.ZN (n_0_180_17), .A (sps__n62));
INV_X1 i_0_180_12 (.ZN (n_0_180_16), .A (sps__n74));
INV_X1 i_0_180_11 (.ZN (n_0_180_15), .A (sps__n86));
NAND4_X1 i_0_180_6 (.ZN (n_0_180_14), .A1 (n_0_180_17), .A2 (n_0_180_16), .A3 (n_0_180_15), .A4 (sps__n2));
INV_X1 i_0_180_5 (.ZN (n_0_180_13), .A (sps__n123));
INV_X1 i_0_180_4 (.ZN (n_0_180_12), .A (sps__n98));
NAND3_X1 i_0_180_1 (.ZN (n_0_180_11), .A1 (n_0_180_13), .A2 (n_0_180_12), .A3 (sps__n112));
INV_X1 i_0_180_0 (.ZN (n_0_180_10), .A (n_0_180_11));
INV_X1 i_0_180_16 (.ZN (n_0_180_9), .A (sps__n68));
INV_X1 i_0_180_15 (.ZN (n_0_180_8), .A (sps__n19));
INV_X1 i_0_180_14 (.ZN (n_0_180_7), .A (address[4]));
INV_X1 i_0_180_13 (.ZN (n_0_180_6), .A (sps__n103));
NAND4_X1 i_0_180_3 (.ZN (n_0_180_5), .A1 (n_0_180_9), .A2 (n_0_180_8), .A3 (n_0_180_7), .A4 (n_0_180_6));
INV_X1 i_0_180_10 (.ZN (n_0_180_4), .A (sps__n55));
INV_X1 i_0_180_9 (.ZN (n_0_180_3), .A (sps__n25));
INV_X1 i_0_180_8 (.ZN (n_0_180_2), .A (sps__n42));
INV_X1 i_0_180_7 (.ZN (n_0_180_1), .A (sps__n92));
NAND4_X1 i_0_180_2 (.ZN (n_0_180_0), .A1 (n_0_180_4), .A2 (n_0_180_3), .A3 (n_0_180_2), .A4 (n_0_180_1));
NAND3_X1 i_0_163_31 (.ZN (n_0_163_30), .A1 (n_0_163_27), .A2 (n_0_163_28), .A3 (n_0_163_29));
NOR2_X1 i_0_163_30 (.ZN (n_0_163_29), .A1 (n_0_163_13), .A2 (n_0_163_23));
NOR2_X1 i_0_163_29 (.ZN (n_0_163_28), .A1 (n_0_163_22), .A2 (n_0_163_21));
NOR2_X1 i_0_163_28 (.ZN (n_0_163_27), .A1 (n_0_163_17), .A2 (n_0_163_20));
NOR2_X1 i_0_163_27 (.ZN (n_0_163_26), .A1 (n_0_163_17), .A2 (n_0_163_13));
NOR2_X1 i_0_163_26 (.ZN (n_0_163_25), .A1 (n_0_163_20), .A2 (n_0_163_21));
NOR2_X1 i_0_163_25 (.ZN (n_0_163_24), .A1 (n_0_163_22), .A2 (n_0_163_23));
NAND3_X1 i_0_163_24 (.ZN (n_0_163_23), .A1 (n_0_163_4), .A2 (n_0_163_2), .A3 (n_0_163_6));
NAND3_X1 i_0_163_23 (.ZN (n_0_163_22), .A1 (n_0_163_1), .A2 (n_0_163_3), .A3 (n_0_163_5));
NAND3_X1 i_0_163_22 (.ZN (n_0_163_21), .A1 (n_0_163_10), .A2 (n_0_163_8), .A3 (n_0_163_12));
NAND3_X1 i_0_163_21 (.ZN (n_0_163_20), .A1 (n_0_163_7), .A2 (n_0_163_9), .A3 (n_0_163_11));
NAND2_X1 i_0_163_20 (.ZN (n_0_163_19), .A1 (n_0_163_30), .A2 (\mem[3][5] ));
INV_X1 i_0_163_19 (.ZN (n_0_163_18), .A (sps__n123));
NAND4_X1 i_0_163_18 (.ZN (n_0_163_17), .A1 (n_0_163_18), .A2 (sps__n2), .A3 (sps__n112), .A4 (sps__n98));
INV_X1 i_0_163_17 (.ZN (n_0_163_16), .A (address[5]));
INV_X1 i_0_163_16 (.ZN (n_0_163_15), .A (address[4]));
INV_X1 i_0_163_15 (.ZN (n_0_163_14), .A (sps__n103));
NAND3_X1 i_0_163_14 (.ZN (n_0_163_13), .A1 (n_0_163_16), .A2 (n_0_163_15), .A3 (n_0_163_14));
INV_X1 i_0_163_13 (.ZN (n_0_163_12), .A (sps__n62));
INV_X1 i_0_163_12 (.ZN (n_0_163_11), .A (sps__n74));
INV_X1 i_0_163_11 (.ZN (n_0_163_10), .A (sps__n7));
INV_X1 i_0_163_10 (.ZN (n_0_163_9), .A (sps__n14));
INV_X1 i_0_163_9 (.ZN (n_0_163_8), .A (sps__n86));
INV_X1 i_0_163_8 (.ZN (n_0_163_7), .A (address[14]));
INV_X1 i_0_163_7 (.ZN (n_0_163_6), .A (sps__n92));
INV_X1 i_0_163_6 (.ZN (n_0_163_5), .A (sps__n68));
INV_X1 i_0_163_5 (.ZN (n_0_163_4), .A (sps__n25));
INV_X1 i_0_163_4 (.ZN (n_0_163_3), .A (sps__n42));
INV_X1 i_0_163_3 (.ZN (n_0_163_2), .A (sps__n51));
INV_X1 i_0_163_2 (.ZN (n_0_163_1), .A (sps__n55));
NAND4_X1 i_0_163_1 (.ZN (n_0_163_0), .A1 (n_0_163_26), .A2 (n_0_163_25), .A3 (n_0_163_24), .A4 (data[5]));
NAND2_X1 i_0_163_0 (.ZN (n_0_154), .A1 (n_0_163_19), .A2 (n_0_163_0));
NAND3_X1 i_0_146_36 (.ZN (n_0_153), .A1 (n_0_146_33), .A2 (n_0_146_34), .A3 (n_0_146_35));
NAND2_X1 i_0_146_35 (.ZN (n_0_146_35), .A1 (n_0_146_24), .A2 (\mem[4][5] ));
NAND2_X1 i_0_146_34 (.ZN (n_0_146_34), .A1 (n_0_146_23), .A2 (\mem[4][5] ));
NAND3_X1 i_0_146_33 (.ZN (n_0_146_33), .A1 (n_0_146_26), .A2 (n_0_146_32), .A3 (n_0_146_29));
NOR2_X1 i_0_146_32 (.ZN (n_0_146_32), .A1 (n_0_146_0), .A2 (n_0_146_18));
INV_X1 i_0_146_31 (.ZN (n_0_146_31), .A (n_0_146_18));
INV_X1 i_0_146_30 (.ZN (n_0_146_30), .A (n_0_146_0));
NOR2_X1 i_0_146_29 (.ZN (n_0_146_29), .A1 (n_0_146_5), .A2 (n_0_146_14));
INV_X1 i_0_146_28 (.ZN (n_0_146_28), .A (n_0_146_14));
INV_X1 i_0_146_27 (.ZN (n_0_146_27), .A (n_0_146_5));
INV_X1 i_0_146_26 (.ZN (n_0_146_26), .A (n_0_146_25));
NAND2_X1 i_0_146_25 (.ZN (n_0_146_25), .A1 (n_0_146_10), .A2 (data[5]));
NAND2_X1 i_0_146_24 (.ZN (n_0_146_24), .A1 (n_0_146_30), .A2 (n_0_146_27));
NAND3_X1 i_0_146_23 (.ZN (n_0_146_23), .A1 (n_0_146_31), .A2 (n_0_146_28), .A3 (n_0_146_10));
INV_X1 i_0_146_22 (.ZN (n_0_146_22), .A (address[14]));
INV_X1 i_0_146_21 (.ZN (n_0_146_21), .A (sps__n9));
INV_X1 i_0_146_20 (.ZN (n_0_146_20), .A (sps__n15));
INV_X1 i_0_146_19 (.ZN (n_0_146_19), .A (sps__n51));
NAND4_X1 i_0_146_18 (.ZN (n_0_146_18), .A1 (n_0_146_22), .A2 (n_0_146_21), .A3 (n_0_146_20), .A4 (n_0_146_19));
INV_X1 i_0_146_17 (.ZN (n_0_146_17), .A (sps__n62));
INV_X1 i_0_146_12 (.ZN (n_0_146_16), .A (sps__n75));
INV_X1 i_0_146_11 (.ZN (n_0_146_15), .A (sps__n86));
NAND4_X1 i_0_146_6 (.ZN (n_0_146_14), .A1 (n_0_146_17), .A2 (n_0_146_16), .A3 (n_0_146_15), .A4 (sps__n2));
INV_X1 i_0_146_5 (.ZN (n_0_146_13), .A (sps__n112));
INV_X1 i_0_146_4 (.ZN (n_0_146_12), .A (sps__n98));
NAND3_X1 i_0_146_1 (.ZN (n_0_146_11), .A1 (n_0_146_13), .A2 (n_0_146_12), .A3 (sps__n123));
INV_X1 i_0_146_0 (.ZN (n_0_146_10), .A (n_0_146_11));
INV_X1 i_0_146_16 (.ZN (n_0_146_9), .A (sps__n68));
INV_X1 i_0_146_15 (.ZN (n_0_146_8), .A (address[5]));
INV_X1 i_0_146_14 (.ZN (n_0_146_7), .A (sps__n81));
INV_X1 i_0_146_13 (.ZN (n_0_146_6), .A (sps__n105));
NAND4_X1 i_0_146_3 (.ZN (n_0_146_5), .A1 (n_0_146_9), .A2 (n_0_146_8), .A3 (n_0_146_7), .A4 (n_0_146_6));
INV_X1 i_0_146_10 (.ZN (n_0_146_4), .A (sps__n55));
INV_X1 i_0_146_9 (.ZN (n_0_146_3), .A (sps__n25));
INV_X1 i_0_146_8 (.ZN (n_0_146_2), .A (sps__n42));
INV_X1 i_0_146_7 (.ZN (n_0_146_1), .A (sps__n92));
NAND4_X1 i_0_146_2 (.ZN (n_0_146_0), .A1 (n_0_146_4), .A2 (n_0_146_3), .A3 (n_0_146_2), .A4 (n_0_146_1));
NAND3_X1 i_0_129_31 (.ZN (n_0_129_30), .A1 (n_0_129_27), .A2 (n_0_129_28), .A3 (n_0_129_29));
NOR2_X1 i_0_129_30 (.ZN (n_0_129_29), .A1 (n_0_129_13), .A2 (n_0_129_23));
NOR2_X1 i_0_129_29 (.ZN (n_0_129_28), .A1 (n_0_129_22), .A2 (n_0_129_21));
NOR2_X1 i_0_129_28 (.ZN (n_0_129_27), .A1 (n_0_129_17), .A2 (n_0_129_20));
NOR2_X1 i_0_129_27 (.ZN (n_0_129_26), .A1 (n_0_129_17), .A2 (n_0_129_13));
NOR2_X1 i_0_129_26 (.ZN (n_0_129_25), .A1 (n_0_129_20), .A2 (n_0_129_21));
NOR2_X1 i_0_129_25 (.ZN (n_0_129_24), .A1 (n_0_129_22), .A2 (n_0_129_23));
NAND3_X1 i_0_129_24 (.ZN (n_0_129_23), .A1 (n_0_129_4), .A2 (n_0_129_2), .A3 (n_0_129_6));
NAND3_X1 i_0_129_23 (.ZN (n_0_129_22), .A1 (n_0_129_1), .A2 (n_0_129_3), .A3 (n_0_129_5));
NAND3_X1 i_0_129_22 (.ZN (n_0_129_21), .A1 (n_0_129_10), .A2 (n_0_129_8), .A3 (n_0_129_12));
NAND3_X1 i_0_129_21 (.ZN (n_0_129_20), .A1 (n_0_129_7), .A2 (n_0_129_9), .A3 (n_0_129_11));
NAND2_X1 i_0_129_20 (.ZN (n_0_129_19), .A1 (n_0_129_30), .A2 (\mem[5][5] ));
INV_X1 i_0_129_19 (.ZN (n_0_129_18), .A (sps__n112));
NAND4_X1 i_0_129_18 (.ZN (n_0_129_17), .A1 (n_0_129_18), .A2 (sps__n2), .A3 (sps__n123), .A4 (sps__n98));
INV_X1 i_0_129_17 (.ZN (n_0_129_16), .A (address[5]));
INV_X1 i_0_129_16 (.ZN (n_0_129_15), .A (address[4]));
INV_X1 i_0_129_15 (.ZN (n_0_129_14), .A (sps__n103));
NAND3_X1 i_0_129_14 (.ZN (n_0_129_13), .A1 (n_0_129_16), .A2 (n_0_129_15), .A3 (n_0_129_14));
INV_X1 i_0_129_13 (.ZN (n_0_129_12), .A (sps__n62));
INV_X1 i_0_129_12 (.ZN (n_0_129_11), .A (sps__n74));
INV_X1 i_0_129_11 (.ZN (n_0_129_10), .A (sps__n7));
INV_X1 i_0_129_10 (.ZN (n_0_129_9), .A (sps__n15));
INV_X1 i_0_129_9 (.ZN (n_0_129_8), .A (sps__n86));
INV_X1 i_0_129_8 (.ZN (n_0_129_7), .A (address[14]));
INV_X1 i_0_129_7 (.ZN (n_0_129_6), .A (sps__n92));
INV_X1 i_0_129_6 (.ZN (n_0_129_5), .A (sps__n68));
INV_X1 i_0_129_5 (.ZN (n_0_129_4), .A (sps__n25));
INV_X1 i_0_129_4 (.ZN (n_0_129_3), .A (sps__n42));
INV_X1 i_0_129_3 (.ZN (n_0_129_2), .A (sps__n51));
INV_X1 i_0_129_2 (.ZN (n_0_129_1), .A (sps__n55));
NAND4_X1 i_0_129_1 (.ZN (n_0_129_0), .A1 (n_0_129_26), .A2 (n_0_129_25), .A3 (n_0_129_24), .A4 (data[5]));
NAND2_X1 i_0_129_0 (.ZN (n_0_152), .A1 (n_0_129_19), .A2 (n_0_129_0));
NAND3_X1 i_0_112_31 (.ZN (n_0_112_30), .A1 (n_0_112_27), .A2 (n_0_112_28), .A3 (n_0_112_29));
NOR2_X1 i_0_112_30 (.ZN (n_0_112_29), .A1 (n_0_112_13), .A2 (n_0_112_23));
NOR2_X1 i_0_112_29 (.ZN (n_0_112_28), .A1 (n_0_112_22), .A2 (n_0_112_21));
NOR2_X1 i_0_112_28 (.ZN (n_0_112_27), .A1 (n_0_112_17), .A2 (n_0_112_20));
NOR2_X1 i_0_112_27 (.ZN (n_0_112_26), .A1 (n_0_112_17), .A2 (n_0_112_13));
NOR2_X1 i_0_112_26 (.ZN (n_0_112_25), .A1 (n_0_112_20), .A2 (n_0_112_21));
NOR2_X1 i_0_112_25 (.ZN (n_0_112_24), .A1 (n_0_112_22), .A2 (n_0_112_23));
NAND3_X1 i_0_112_24 (.ZN (n_0_112_23), .A1 (n_0_112_4), .A2 (n_0_112_2), .A3 (n_0_112_6));
NAND3_X1 i_0_112_23 (.ZN (n_0_112_22), .A1 (n_0_112_1), .A2 (n_0_112_3), .A3 (n_0_112_5));
NAND3_X1 i_0_112_22 (.ZN (n_0_112_21), .A1 (n_0_112_10), .A2 (n_0_112_8), .A3 (n_0_112_12));
NAND3_X1 i_0_112_21 (.ZN (n_0_112_20), .A1 (n_0_112_7), .A2 (n_0_112_9), .A3 (n_0_112_11));
NAND2_X1 i_0_112_20 (.ZN (n_0_112_19), .A1 (n_0_112_30), .A2 (\mem[6][5] ));
INV_X1 i_0_112_19 (.ZN (n_0_112_18), .A (sps__n98));
NAND4_X1 i_0_112_18 (.ZN (n_0_112_17), .A1 (n_0_112_18), .A2 (sps__n2), .A3 (sps__n123), .A4 (sps__n112));
INV_X1 i_0_112_17 (.ZN (n_0_112_16), .A (sps__n19));
INV_X1 i_0_112_16 (.ZN (n_0_112_15), .A (sps__n81));
INV_X1 i_0_112_15 (.ZN (n_0_112_14), .A (sps__n105));
NAND3_X1 i_0_112_14 (.ZN (n_0_112_13), .A1 (n_0_112_16), .A2 (n_0_112_15), .A3 (n_0_112_14));
INV_X1 i_0_112_13 (.ZN (n_0_112_12), .A (sps__n62));
INV_X1 i_0_112_12 (.ZN (n_0_112_11), .A (sps__n75));
INV_X1 i_0_112_11 (.ZN (n_0_112_10), .A (sps__n9));
INV_X1 i_0_112_10 (.ZN (n_0_112_9), .A (sps__n15));
INV_X1 i_0_112_9 (.ZN (n_0_112_8), .A (sps__n86));
INV_X1 i_0_112_8 (.ZN (n_0_112_7), .A (address[14]));
INV_X1 i_0_112_7 (.ZN (n_0_112_6), .A (sps__n92));
INV_X1 i_0_112_6 (.ZN (n_0_112_5), .A (sps__n68));
INV_X1 i_0_112_5 (.ZN (n_0_112_4), .A (sps__n28));
INV_X1 i_0_112_4 (.ZN (n_0_112_3), .A (sps__n42));
INV_X1 i_0_112_3 (.ZN (n_0_112_2), .A (sps__n51));
INV_X1 i_0_112_2 (.ZN (n_0_112_1), .A (sps__n55));
NAND4_X1 i_0_112_1 (.ZN (n_0_112_0), .A1 (n_0_112_26), .A2 (n_0_112_25), .A3 (n_0_112_24), .A4 (data[5]));
NAND2_X1 i_0_112_0 (.ZN (n_0_149), .A1 (n_0_112_19), .A2 (n_0_112_0));
NAND3_X1 i_0_95_27 (.ZN (n_0_95_26), .A1 (n_0_95_23), .A2 (n_0_95_24), .A3 (n_0_95_25));
NOR2_X1 i_0_95_26 (.ZN (n_0_95_25), .A1 (n_0_95_17), .A2 (n_0_95_13));
NOR2_X1 i_0_95_25 (.ZN (n_0_95_24), .A1 (n_0_95_19), .A2 (n_0_95_20));
NOR2_X1 i_0_95_24 (.ZN (n_0_95_23), .A1 (n_0_95_21), .A2 (n_0_95_22));
NAND3_X1 i_0_95_23 (.ZN (n_0_95_22), .A1 (n_0_95_4), .A2 (n_0_95_2), .A3 (n_0_95_6));
NAND3_X1 i_0_95_22 (.ZN (n_0_95_21), .A1 (n_0_95_1), .A2 (n_0_95_3), .A3 (n_0_95_5));
NAND3_X1 i_0_95_21 (.ZN (n_0_95_20), .A1 (n_0_95_10), .A2 (n_0_95_8), .A3 (n_0_95_12));
NAND3_X1 i_0_95_20 (.ZN (n_0_95_19), .A1 (n_0_95_7), .A2 (n_0_95_9), .A3 (n_0_95_11));
NAND2_X1 i_0_95_19 (.ZN (n_0_95_18), .A1 (n_0_95_26), .A2 (\mem[7][5] ));
NAND4_X1 i_0_95_18 (.ZN (n_0_95_17), .A1 (sps__n2), .A2 (sps__n123), .A3 (sps__n112), .A4 (sps__n98));
INV_X1 i_0_95_17 (.ZN (n_0_95_16), .A (address[5]));
INV_X1 i_0_95_16 (.ZN (n_0_95_15), .A (address[4]));
INV_X1 i_0_95_15 (.ZN (n_0_95_14), .A (sps__n103));
NAND3_X1 i_0_95_14 (.ZN (n_0_95_13), .A1 (n_0_95_16), .A2 (n_0_95_15), .A3 (n_0_95_14));
INV_X1 i_0_95_13 (.ZN (n_0_95_12), .A (sps__n62));
INV_X1 i_0_95_12 (.ZN (n_0_95_11), .A (sps__n74));
INV_X1 i_0_95_11 (.ZN (n_0_95_10), .A (sps__n7));
INV_X1 i_0_95_10 (.ZN (n_0_95_9), .A (sps__n14));
INV_X1 i_0_95_9 (.ZN (n_0_95_8), .A (sps__n86));
INV_X1 i_0_95_8 (.ZN (n_0_95_7), .A (address[14]));
INV_X1 i_0_95_7 (.ZN (n_0_95_6), .A (sps__n92));
INV_X1 i_0_95_6 (.ZN (n_0_95_5), .A (sps__n68));
INV_X1 i_0_95_5 (.ZN (n_0_95_4), .A (address[9]));
INV_X1 i_0_95_4 (.ZN (n_0_95_3), .A (sps__n42));
INV_X1 i_0_95_3 (.ZN (n_0_95_2), .A (sps__n51));
INV_X1 i_0_95_2 (.ZN (n_0_95_1), .A (sps__n55));
NAND4_X1 i_0_95_1 (.ZN (n_0_95_0), .A1 (n_0_95_25), .A2 (n_0_95_24), .A3 (n_0_95_23), .A4 (data[5]));
NAND2_X1 i_0_95_0 (.ZN (n_0_148), .A1 (n_0_95_18), .A2 (n_0_95_0));
NAND3_X1 i_0_78_35 (.ZN (n_0_147), .A1 (n_0_78_32), .A2 (n_0_78_33), .A3 (n_0_78_34));
NAND2_X1 i_0_78_34 (.ZN (n_0_78_34), .A1 (n_0_78_23), .A2 (\mem[8][5] ));
NAND3_X1 i_0_78_29 (.ZN (n_0_78_33), .A1 (n_0_78_26), .A2 (n_0_78_31), .A3 (n_0_78_28));
NAND2_X1 i_0_78_28 (.ZN (n_0_78_32), .A1 (n_0_78_27), .A2 (\mem[8][5] ));
NOR2_X1 i_0_78_24 (.ZN (n_0_78_31), .A1 (n_0_78_18), .A2 (n_0_78_0));
INV_X1 i_0_78_23 (.ZN (n_0_78_30), .A (n_0_78_0));
INV_X1 i_0_78_22 (.ZN (n_0_78_29), .A (n_0_78_18));
INV_X1 i_0_78_21 (.ZN (n_0_78_28), .A (n_0_78_5));
NAND3_X1 i_0_78_20 (.ZN (n_0_78_27), .A1 (n_0_78_28), .A2 (n_0_78_30), .A3 (n_0_78_9));
NOR2_X1 i_0_78_19 (.ZN (n_0_78_26), .A1 (n_0_78_14), .A2 (n_0_78_24));
INV_X1 i_0_78_18 (.ZN (n_0_78_25), .A (n_0_78_14));
NAND2_X1 i_0_78_17 (.ZN (n_0_78_24), .A1 (n_0_78_9), .A2 (data[5]));
NAND2_X1 i_0_78_16 (.ZN (n_0_78_23), .A1 (n_0_78_29), .A2 (n_0_78_25));
INV_X1 i_0_78_33 (.ZN (n_0_78_22), .A (address[14]));
INV_X1 i_0_78_32 (.ZN (n_0_78_21), .A (sps__n7));
INV_X1 i_0_78_31 (.ZN (n_0_78_20), .A (sps__n15));
INV_X1 i_0_78_30 (.ZN (n_0_78_19), .A (sps__n51));
NAND4_X1 i_0_78_3 (.ZN (n_0_78_18), .A1 (n_0_78_22), .A2 (n_0_78_21), .A3 (n_0_78_20), .A4 (n_0_78_19));
INV_X1 i_0_78_27 (.ZN (n_0_78_17), .A (sps__n62));
INV_X1 i_0_78_26 (.ZN (n_0_78_16), .A (sps__n75));
INV_X1 i_0_78_25 (.ZN (n_0_78_15), .A (sps__n86));
NAND4_X1 i_0_78_8 (.ZN (n_0_78_14), .A1 (n_0_78_17), .A2 (n_0_78_16), .A3 (n_0_78_15), .A4 (sps__n2));
INV_X1 i_0_78_15 (.ZN (n_0_78_13), .A (sps__n123));
INV_X1 i_0_78_14 (.ZN (n_0_78_12), .A (sps__n112));
INV_X1 i_0_78_13 (.ZN (n_0_78_11), .A (sps__n98));
NAND3_X1 i_0_78_12 (.ZN (n_0_78_10), .A1 (n_0_78_13), .A2 (n_0_78_12), .A3 (n_0_78_11));
INV_X1 i_0_78_11 (.ZN (n_0_78_9), .A (n_0_78_10));
INV_X1 i_0_78_10 (.ZN (n_0_78_8), .A (sps__n68));
INV_X1 i_0_78_9 (.ZN (n_0_78_7), .A (address[5]));
INV_X1 i_0_78_7 (.ZN (n_0_78_6), .A (sps__n81));
NAND4_X1 i_0_78_6 (.ZN (n_0_78_5), .A1 (n_0_78_8), .A2 (n_0_78_7), .A3 (n_0_78_6), .A4 (sps__n105));
INV_X1 i_0_78_5 (.ZN (n_0_78_4), .A (sps__n55));
INV_X1 i_0_78_4 (.ZN (n_0_78_3), .A (sps__n25));
INV_X1 i_0_78_2 (.ZN (n_0_78_2), .A (sps__n42));
INV_X1 i_0_78_1 (.ZN (n_0_78_1), .A (sps__n92));
NAND4_X1 i_0_78_0 (.ZN (n_0_78_0), .A1 (n_0_78_4), .A2 (n_0_78_3), .A3 (n_0_78_2), .A4 (n_0_78_1));
NOR2_X1 i_0_61_34 (.ZN (n_0_61_33), .A1 (n_0_61_19), .A2 (n_0_61_0));
INV_X1 i_0_61_33 (.ZN (n_0_61_32), .A (n_0_61_0));
INV_X1 i_0_61_28 (.ZN (n_0_61_31), .A (n_0_61_19));
NAND2_X1 i_0_61_27 (.ZN (n_0_61_30), .A1 (n_0_61_29), .A2 (\mem[9][5] ));
NAND3_X1 i_0_61_23 (.ZN (n_0_61_29), .A1 (n_0_61_5), .A2 (n_0_61_32), .A3 (n_0_61_10));
NAND3_X1 i_0_61_22 (.ZN (n_0_61_28), .A1 (n_0_61_27), .A2 (n_0_61_33), .A3 (n_0_61_14));
NOR2_X1 i_0_61_21 (.ZN (n_0_61_27), .A1 (n_0_61_6), .A2 (n_0_61_26));
NAND2_X1 i_0_61_20 (.ZN (n_0_61_26), .A1 (n_0_61_10), .A2 (data[5]));
NAND2_X1 i_0_61_19 (.ZN (n_0_61_25), .A1 (n_0_61_31), .A2 (n_0_61_14));
NAND3_X1 i_0_61_18 (.ZN (n_0_146), .A1 (n_0_61_28), .A2 (n_0_61_30), .A3 (n_0_61_24));
NAND2_X1 i_0_61_17 (.ZN (n_0_61_24), .A1 (n_0_61_25), .A2 (\mem[9][5] ));
INV_X1 i_0_61_32 (.ZN (n_0_61_23), .A (address[14]));
INV_X1 i_0_61_31 (.ZN (n_0_61_22), .A (sps__n7));
INV_X1 i_0_61_30 (.ZN (n_0_61_21), .A (sps__n14));
INV_X1 i_0_61_29 (.ZN (n_0_61_20), .A (sps__n51));
NAND4_X1 i_0_61_3 (.ZN (n_0_61_19), .A1 (n_0_61_23), .A2 (n_0_61_22), .A3 (n_0_61_21), .A4 (n_0_61_20));
INV_X1 i_0_61_26 (.ZN (n_0_61_18), .A (sps__n62));
INV_X1 i_0_61_25 (.ZN (n_0_61_17), .A (sps__n74));
INV_X1 i_0_61_24 (.ZN (n_0_61_16), .A (sps__n86));
NAND4_X1 i_0_61_6 (.ZN (n_0_61_15), .A1 (n_0_61_18), .A2 (n_0_61_17), .A3 (n_0_61_16), .A4 (sps__n2));
INV_X1 i_0_61_16 (.ZN (n_0_61_14), .A (n_0_61_15));
INV_X1 i_0_61_15 (.ZN (n_0_61_13), .A (sps__n123));
INV_X1 i_0_61_14 (.ZN (n_0_61_12), .A (sps__n114));
NAND3_X1 i_0_61_13 (.ZN (n_0_61_11), .A1 (n_0_61_13), .A2 (n_0_61_12), .A3 (sps__n98));
INV_X1 i_0_61_12 (.ZN (n_0_61_10), .A (n_0_61_11));
INV_X1 i_0_61_11 (.ZN (n_0_61_9), .A (sps__n68));
INV_X1 i_0_61_10 (.ZN (n_0_61_8), .A (address[5]));
INV_X1 i_0_61_9 (.ZN (n_0_61_7), .A (address[4]));
NAND4_X1 i_0_61_8 (.ZN (n_0_61_6), .A1 (n_0_61_9), .A2 (n_0_61_8), .A3 (n_0_61_7), .A4 (sps__n103));
INV_X1 i_0_61_7 (.ZN (n_0_61_5), .A (n_0_61_6));
INV_X1 i_0_61_5 (.ZN (n_0_61_4), .A (sps__n55));
INV_X1 i_0_61_4 (.ZN (n_0_61_3), .A (address[9]));
INV_X1 i_0_61_2 (.ZN (n_0_61_2), .A (sps__n42));
INV_X1 i_0_61_1 (.ZN (n_0_61_1), .A (sps__n92));
NAND4_X1 i_0_61_0 (.ZN (n_0_61_0), .A1 (n_0_61_4), .A2 (n_0_61_3), .A3 (n_0_61_2), .A4 (n_0_61_1));
NOR2_X1 i_0_44_34 (.ZN (n_0_44_33), .A1 (n_0_44_19), .A2 (n_0_44_0));
INV_X1 i_0_44_33 (.ZN (n_0_44_32), .A (n_0_44_0));
INV_X1 i_0_44_28 (.ZN (n_0_44_31), .A (n_0_44_19));
NAND2_X1 i_0_44_27 (.ZN (n_0_44_30), .A1 (n_0_44_29), .A2 (\mem[10][5] ));
NAND3_X1 i_0_44_23 (.ZN (n_0_44_29), .A1 (n_0_44_5), .A2 (n_0_44_32), .A3 (n_0_44_10));
NAND3_X1 i_0_44_22 (.ZN (n_0_44_28), .A1 (n_0_44_27), .A2 (n_0_44_33), .A3 (n_0_44_14));
NOR2_X1 i_0_44_21 (.ZN (n_0_44_27), .A1 (n_0_44_6), .A2 (n_0_44_26));
NAND2_X1 i_0_44_20 (.ZN (n_0_44_26), .A1 (n_0_44_10), .A2 (data[5]));
NAND2_X1 i_0_44_19 (.ZN (n_0_44_25), .A1 (n_0_44_31), .A2 (n_0_44_14));
NAND3_X1 i_0_44_18 (.ZN (n_0_145), .A1 (n_0_44_28), .A2 (n_0_44_30), .A3 (n_0_44_24));
NAND2_X1 i_0_44_17 (.ZN (n_0_44_24), .A1 (n_0_44_25), .A2 (\mem[10][5] ));
INV_X1 i_0_44_32 (.ZN (n_0_44_23), .A (address[14]));
INV_X1 i_0_44_31 (.ZN (n_0_44_22), .A (sps__n9));
INV_X1 i_0_44_30 (.ZN (n_0_44_21), .A (sps__n15));
INV_X1 i_0_44_29 (.ZN (n_0_44_20), .A (sps__n51));
NAND4_X1 i_0_44_3 (.ZN (n_0_44_19), .A1 (n_0_44_23), .A2 (n_0_44_22), .A3 (n_0_44_21), .A4 (n_0_44_20));
INV_X1 i_0_44_26 (.ZN (n_0_44_18), .A (sps__n62));
INV_X1 i_0_44_25 (.ZN (n_0_44_17), .A (sps__n75));
INV_X1 i_0_44_24 (.ZN (n_0_44_16), .A (sps__n86));
NAND4_X1 i_0_44_6 (.ZN (n_0_44_15), .A1 (n_0_44_18), .A2 (n_0_44_17), .A3 (n_0_44_16), .A4 (sps__n2));
INV_X1 i_0_44_16 (.ZN (n_0_44_14), .A (n_0_44_15));
INV_X1 i_0_44_15 (.ZN (n_0_44_13), .A (sps__n123));
INV_X1 i_0_44_14 (.ZN (n_0_44_12), .A (sps__n98));
NAND3_X1 i_0_44_13 (.ZN (n_0_44_11), .A1 (n_0_44_13), .A2 (n_0_44_12), .A3 (sps__n112));
INV_X1 i_0_44_12 (.ZN (n_0_44_10), .A (n_0_44_11));
INV_X1 i_0_44_11 (.ZN (n_0_44_9), .A (sps__n68));
INV_X1 i_0_44_10 (.ZN (n_0_44_8), .A (sps__n19));
INV_X1 i_0_44_9 (.ZN (n_0_44_7), .A (sps__n81));
NAND4_X1 i_0_44_8 (.ZN (n_0_44_6), .A1 (n_0_44_9), .A2 (n_0_44_8), .A3 (n_0_44_7), .A4 (sps__n105));
INV_X1 i_0_44_7 (.ZN (n_0_44_5), .A (n_0_44_6));
INV_X1 i_0_44_5 (.ZN (n_0_44_4), .A (sps__n55));
INV_X1 i_0_44_4 (.ZN (n_0_44_3), .A (sps__n28));
INV_X1 i_0_44_2 (.ZN (n_0_44_2), .A (sps__n43));
INV_X1 i_0_44_1 (.ZN (n_0_44_1), .A (sps__n92));
NAND4_X1 i_0_44_0 (.ZN (n_0_44_0), .A1 (n_0_44_4), .A2 (n_0_44_3), .A3 (n_0_44_2), .A4 (n_0_44_1));
NAND3_X1 i_0_27_37 (.ZN (n_0_144), .A1 (n_0_27_34), .A2 (n_0_27_35), .A3 (n_0_27_36));
NAND2_X1 i_0_27_36 (.ZN (n_0_27_36), .A1 (n_0_27_25), .A2 (\mem[0][6] ));
NAND3_X1 i_0_27_35 (.ZN (n_0_27_35), .A1 (n_0_27_27), .A2 (n_0_27_33), .A3 (n_0_27_30));
NAND2_X1 i_0_27_34 (.ZN (n_0_27_34), .A1 (n_0_27_24), .A2 (\mem[0][6] ));
NOR2_X1 i_0_27_33 (.ZN (n_0_27_33), .A1 (n_0_27_0), .A2 (n_0_27_19));
INV_X1 i_0_27_32 (.ZN (n_0_27_32), .A (n_0_27_19));
INV_X1 i_0_27_31 (.ZN (n_0_27_31), .A (n_0_27_0));
NOR2_X1 i_0_27_30 (.ZN (n_0_27_30), .A1 (n_0_27_5), .A2 (n_0_27_15));
INV_X1 i_0_27_29 (.ZN (n_0_27_29), .A (n_0_27_15));
INV_X1 i_0_27_28 (.ZN (n_0_27_28), .A (n_0_27_5));
INV_X1 i_0_27_27 (.ZN (n_0_27_27), .A (n_0_27_26));
NAND2_X1 i_0_27_26 (.ZN (n_0_27_26), .A1 (n_0_27_10), .A2 (data[6]));
NAND2_X1 i_0_27_25 (.ZN (n_0_27_25), .A1 (n_0_27_31), .A2 (n_0_27_28));
NAND3_X1 i_0_27_24 (.ZN (n_0_27_24), .A1 (n_0_27_32), .A2 (n_0_27_29), .A3 (n_0_27_10));
INV_X1 i_0_27_23 (.ZN (n_0_27_23), .A (sps__n36));
INV_X1 i_0_27_22 (.ZN (n_0_27_22), .A (sps__n7));
INV_X1 i_0_27_21 (.ZN (n_0_27_21), .A (sps__n13));
INV_X1 i_0_27_20 (.ZN (n_0_27_20), .A (address[11]));
NAND4_X1 i_0_27_19 (.ZN (n_0_27_19), .A1 (n_0_27_23), .A2 (n_0_27_22), .A3 (n_0_27_21), .A4 (n_0_27_20));
INV_X1 i_0_27_18 (.ZN (n_0_27_18), .A (sps__n61));
INV_X1 i_0_27_17 (.ZN (n_0_27_17), .A (sps__n73));
INV_X1 i_0_27_12 (.ZN (n_0_27_16), .A (sps__n85));
NAND4_X1 i_0_27_11 (.ZN (n_0_27_15), .A1 (n_0_27_18), .A2 (n_0_27_17), .A3 (n_0_27_16), .A4 (sps__n1));
INV_X1 i_0_27_6 (.ZN (n_0_27_14), .A (address[2]));
INV_X1 i_0_27_5 (.ZN (n_0_27_13), .A (sps__n113));
INV_X1 i_0_27_4 (.ZN (n_0_27_12), .A (sps__n97));
NAND3_X1 i_0_27_1 (.ZN (n_0_27_11), .A1 (n_0_27_14), .A2 (n_0_27_13), .A3 (n_0_27_12));
INV_X1 i_0_27_0 (.ZN (n_0_27_10), .A (n_0_27_11));
INV_X1 i_0_27_16 (.ZN (n_0_27_9), .A (sps__n69));
INV_X1 i_0_27_15 (.ZN (n_0_27_8), .A (sps__n20));
INV_X1 i_0_27_14 (.ZN (n_0_27_7), .A (sps__n79));
INV_X1 i_0_27_13 (.ZN (n_0_27_6), .A (sps__n106));
NAND4_X1 i_0_27_3 (.ZN (n_0_27_5), .A1 (n_0_27_9), .A2 (n_0_27_8), .A3 (n_0_27_7), .A4 (n_0_27_6));
INV_X1 i_0_27_10 (.ZN (n_0_27_4), .A (sps__n56));
INV_X1 i_0_27_9 (.ZN (n_0_27_3), .A (sps__n27));
INV_X1 i_0_27_8 (.ZN (n_0_27_2), .A (sps__n41));
INV_X1 i_0_27_7 (.ZN (n_0_27_1), .A (sps__n93));
NAND4_X1 i_0_27_2 (.ZN (n_0_27_0), .A1 (n_0_27_4), .A2 (n_0_27_3), .A3 (n_0_27_2), .A4 (n_0_27_1));
NAND3_X1 i_0_42_36 (.ZN (n_0_143), .A1 (n_0_42_33), .A2 (n_0_42_34), .A3 (n_0_42_35));
NAND2_X1 i_0_42_35 (.ZN (n_0_42_35), .A1 (n_0_42_24), .A2 (\mem[1][6] ));
NAND2_X1 i_0_42_34 (.ZN (n_0_42_34), .A1 (n_0_42_23), .A2 (\mem[1][6] ));
NAND3_X1 i_0_42_33 (.ZN (n_0_42_33), .A1 (n_0_42_26), .A2 (n_0_42_32), .A3 (n_0_42_29));
NOR2_X1 i_0_42_32 (.ZN (n_0_42_32), .A1 (n_0_42_0), .A2 (n_0_42_18));
INV_X1 i_0_42_31 (.ZN (n_0_42_31), .A (n_0_42_18));
INV_X1 i_0_42_30 (.ZN (n_0_42_30), .A (n_0_42_0));
NOR2_X1 i_0_42_29 (.ZN (n_0_42_29), .A1 (n_0_42_5), .A2 (n_0_42_14));
INV_X1 i_0_42_28 (.ZN (n_0_42_28), .A (n_0_42_14));
INV_X1 i_0_42_27 (.ZN (n_0_42_27), .A (n_0_42_5));
INV_X1 i_0_42_26 (.ZN (n_0_42_26), .A (n_0_42_25));
NAND2_X1 i_0_42_25 (.ZN (n_0_42_25), .A1 (n_0_42_10), .A2 (data[6]));
NAND2_X1 i_0_42_24 (.ZN (n_0_42_24), .A1 (n_0_42_30), .A2 (n_0_42_27));
NAND3_X1 i_0_42_23 (.ZN (n_0_42_23), .A1 (n_0_42_31), .A2 (n_0_42_28), .A3 (n_0_42_10));
INV_X1 i_0_42_22 (.ZN (n_0_42_22), .A (sps__n36));
INV_X1 i_0_42_21 (.ZN (n_0_42_21), .A (sps__n7));
INV_X1 i_0_42_20 (.ZN (n_0_42_20), .A (address[12]));
INV_X1 i_0_42_19 (.ZN (n_0_42_19), .A (address[11]));
NAND4_X1 i_0_42_18 (.ZN (n_0_42_18), .A1 (n_0_42_22), .A2 (n_0_42_21), .A3 (n_0_42_20), .A4 (n_0_42_19));
INV_X1 i_0_42_17 (.ZN (n_0_42_17), .A (RST));
INV_X1 i_0_42_12 (.ZN (n_0_42_16), .A (sps__n73));
INV_X1 i_0_42_11 (.ZN (n_0_42_15), .A (sps__n85));
NAND4_X1 i_0_42_6 (.ZN (n_0_42_14), .A1 (n_0_42_17), .A2 (n_0_42_16), .A3 (n_0_42_15), .A4 (sps__n1));
INV_X1 i_0_42_5 (.ZN (n_0_42_13), .A (sps__n123));
INV_X1 i_0_42_4 (.ZN (n_0_42_12), .A (sps__n114));
NAND3_X1 i_0_42_1 (.ZN (n_0_42_11), .A1 (n_0_42_13), .A2 (n_0_42_12), .A3 (sps__n97));
INV_X1 i_0_42_0 (.ZN (n_0_42_10), .A (n_0_42_11));
INV_X1 i_0_42_16 (.ZN (n_0_42_9), .A (sps__n69));
INV_X1 i_0_42_15 (.ZN (n_0_42_8), .A (sps__n20));
INV_X1 i_0_42_14 (.ZN (n_0_42_7), .A (sps__n79));
INV_X1 i_0_42_13 (.ZN (n_0_42_6), .A (address[3]));
NAND4_X1 i_0_42_3 (.ZN (n_0_42_5), .A1 (n_0_42_9), .A2 (n_0_42_8), .A3 (n_0_42_7), .A4 (n_0_42_6));
INV_X1 i_0_42_10 (.ZN (n_0_42_4), .A (sps__n56));
INV_X1 i_0_42_9 (.ZN (n_0_42_3), .A (sps__n26));
INV_X1 i_0_42_8 (.ZN (n_0_42_2), .A (address[8]));
INV_X1 i_0_42_7 (.ZN (n_0_42_1), .A (address[7]));
NAND4_X1 i_0_42_2 (.ZN (n_0_42_0), .A1 (n_0_42_4), .A2 (n_0_42_3), .A3 (n_0_42_2), .A4 (n_0_42_1));
NAND3_X1 i_0_179_36 (.ZN (n_0_142), .A1 (n_0_179_33), .A2 (n_0_179_34), .A3 (n_0_179_35));
NAND2_X1 i_0_179_35 (.ZN (n_0_179_35), .A1 (n_0_179_24), .A2 (\mem[2][6] ));
NAND2_X1 i_0_179_34 (.ZN (n_0_179_34), .A1 (n_0_179_23), .A2 (\mem[2][6] ));
NAND3_X1 i_0_179_33 (.ZN (n_0_179_33), .A1 (n_0_179_26), .A2 (n_0_179_32), .A3 (n_0_179_29));
NOR2_X1 i_0_179_32 (.ZN (n_0_179_32), .A1 (n_0_179_0), .A2 (n_0_179_18));
INV_X1 i_0_179_31 (.ZN (n_0_179_31), .A (n_0_179_18));
INV_X1 i_0_179_30 (.ZN (n_0_179_30), .A (n_0_179_0));
NOR2_X1 i_0_179_29 (.ZN (n_0_179_29), .A1 (n_0_179_5), .A2 (n_0_179_14));
INV_X1 i_0_179_28 (.ZN (n_0_179_28), .A (n_0_179_14));
INV_X1 i_0_179_27 (.ZN (n_0_179_27), .A (n_0_179_5));
INV_X1 i_0_179_26 (.ZN (n_0_179_26), .A (n_0_179_25));
NAND2_X1 i_0_179_25 (.ZN (n_0_179_25), .A1 (n_0_179_10), .A2 (data[6]));
NAND2_X1 i_0_179_24 (.ZN (n_0_179_24), .A1 (n_0_179_30), .A2 (n_0_179_27));
NAND3_X1 i_0_179_23 (.ZN (n_0_179_23), .A1 (n_0_179_31), .A2 (n_0_179_28), .A3 (n_0_179_10));
INV_X1 i_0_179_22 (.ZN (n_0_179_22), .A (sps__n36));
INV_X1 i_0_179_21 (.ZN (n_0_179_21), .A (sps__n7));
INV_X1 i_0_179_20 (.ZN (n_0_179_20), .A (sps__n13));
INV_X1 i_0_179_19 (.ZN (n_0_179_19), .A (address[11]));
NAND4_X1 i_0_179_18 (.ZN (n_0_179_18), .A1 (n_0_179_22), .A2 (n_0_179_21), .A3 (n_0_179_20), .A4 (n_0_179_19));
INV_X1 i_0_179_17 (.ZN (n_0_179_17), .A (RST));
INV_X1 i_0_179_12 (.ZN (n_0_179_16), .A (read_signal));
INV_X1 i_0_179_11 (.ZN (n_0_179_15), .A (address[15]));
NAND4_X1 i_0_179_6 (.ZN (n_0_179_14), .A1 (n_0_179_17), .A2 (n_0_179_16), .A3 (n_0_179_15), .A4 (sps__n1));
INV_X1 i_0_179_5 (.ZN (n_0_179_13), .A (address[2]));
INV_X1 i_0_179_4 (.ZN (n_0_179_12), .A (sps__n97));
NAND3_X1 i_0_179_1 (.ZN (n_0_179_11), .A1 (n_0_179_13), .A2 (n_0_179_12), .A3 (sps__n113));
INV_X1 i_0_179_0 (.ZN (n_0_179_10), .A (n_0_179_11));
INV_X1 i_0_179_16 (.ZN (n_0_179_9), .A (sps__n69));
INV_X1 i_0_179_15 (.ZN (n_0_179_8), .A (sps__n20));
INV_X1 i_0_179_14 (.ZN (n_0_179_7), .A (sps__n79));
INV_X1 i_0_179_13 (.ZN (n_0_179_6), .A (sps__n106));
NAND4_X1 i_0_179_3 (.ZN (n_0_179_5), .A1 (n_0_179_9), .A2 (n_0_179_8), .A3 (n_0_179_7), .A4 (n_0_179_6));
INV_X1 i_0_179_10 (.ZN (n_0_179_4), .A (sps__n56));
INV_X1 i_0_179_9 (.ZN (n_0_179_3), .A (sps__n27));
INV_X1 i_0_179_8 (.ZN (n_0_179_2), .A (sps__n41));
INV_X1 i_0_179_7 (.ZN (n_0_179_1), .A (sps__n93));
NAND4_X1 i_0_179_2 (.ZN (n_0_179_0), .A1 (n_0_179_4), .A2 (n_0_179_3), .A3 (n_0_179_2), .A4 (n_0_179_1));
NAND3_X1 i_0_162_31 (.ZN (n_0_162_30), .A1 (n_0_162_27), .A2 (n_0_162_28), .A3 (n_0_162_29));
NOR2_X1 i_0_162_30 (.ZN (n_0_162_29), .A1 (n_0_162_13), .A2 (n_0_162_23));
NOR2_X1 i_0_162_29 (.ZN (n_0_162_28), .A1 (n_0_162_22), .A2 (n_0_162_21));
NOR2_X1 i_0_162_28 (.ZN (n_0_162_27), .A1 (n_0_162_17), .A2 (n_0_162_20));
NOR2_X1 i_0_162_27 (.ZN (n_0_162_26), .A1 (n_0_162_17), .A2 (n_0_162_13));
NOR2_X1 i_0_162_26 (.ZN (n_0_162_25), .A1 (n_0_162_20), .A2 (n_0_162_21));
NOR2_X1 i_0_162_25 (.ZN (n_0_162_24), .A1 (n_0_162_22), .A2 (n_0_162_23));
NAND3_X1 i_0_162_24 (.ZN (n_0_162_23), .A1 (n_0_162_4), .A2 (n_0_162_2), .A3 (n_0_162_6));
NAND3_X1 i_0_162_23 (.ZN (n_0_162_22), .A1 (n_0_162_1), .A2 (n_0_162_3), .A3 (n_0_162_5));
NAND3_X1 i_0_162_22 (.ZN (n_0_162_21), .A1 (n_0_162_10), .A2 (n_0_162_8), .A3 (n_0_162_12));
NAND3_X1 i_0_162_21 (.ZN (n_0_162_20), .A1 (n_0_162_7), .A2 (n_0_162_9), .A3 (n_0_162_11));
NAND2_X1 i_0_162_20 (.ZN (n_0_162_19), .A1 (n_0_162_30), .A2 (\mem[3][6] ));
INV_X1 i_0_162_19 (.ZN (n_0_162_18), .A (address[2]));
NAND4_X1 i_0_162_18 (.ZN (n_0_162_17), .A1 (n_0_162_18), .A2 (sps__n1), .A3 (sps__n114), .A4 (sps__n97));
INV_X1 i_0_162_17 (.ZN (n_0_162_16), .A (sps__n20));
INV_X1 i_0_162_16 (.ZN (n_0_162_15), .A (sps__n79));
INV_X1 i_0_162_15 (.ZN (n_0_162_14), .A (address[3]));
NAND3_X1 i_0_162_14 (.ZN (n_0_162_13), .A1 (n_0_162_16), .A2 (n_0_162_15), .A3 (n_0_162_14));
INV_X1 i_0_162_13 (.ZN (n_0_162_12), .A (RST));
INV_X1 i_0_162_12 (.ZN (n_0_162_11), .A (read_signal));
INV_X1 i_0_162_11 (.ZN (n_0_162_10), .A (sps__n7));
INV_X1 i_0_162_10 (.ZN (n_0_162_9), .A (sps__n13));
INV_X1 i_0_162_9 (.ZN (n_0_162_8), .A (sps__n85));
INV_X1 i_0_162_8 (.ZN (n_0_162_7), .A (sps__n36));
INV_X1 i_0_162_7 (.ZN (n_0_162_6), .A (address[7]));
INV_X1 i_0_162_6 (.ZN (n_0_162_5), .A (sps__n69));
INV_X1 i_0_162_5 (.ZN (n_0_162_4), .A (sps__n26));
INV_X1 i_0_162_4 (.ZN (n_0_162_3), .A (address[8]));
INV_X1 i_0_162_3 (.ZN (n_0_162_2), .A (address[11]));
INV_X1 i_0_162_2 (.ZN (n_0_162_1), .A (sps__n56));
NAND4_X1 i_0_162_1 (.ZN (n_0_162_0), .A1 (n_0_162_26), .A2 (n_0_162_25), .A3 (n_0_162_24), .A4 (data[6]));
NAND2_X1 i_0_162_0 (.ZN (n_0_141), .A1 (n_0_162_19), .A2 (n_0_162_0));
NAND3_X1 i_0_145_36 (.ZN (n_0_140), .A1 (n_0_145_33), .A2 (n_0_145_34), .A3 (n_0_145_35));
NAND2_X1 i_0_145_35 (.ZN (n_0_145_35), .A1 (n_0_145_24), .A2 (\mem[4][6] ));
NAND2_X1 i_0_145_34 (.ZN (n_0_145_34), .A1 (n_0_145_23), .A2 (\mem[4][6] ));
NAND3_X1 i_0_145_33 (.ZN (n_0_145_33), .A1 (n_0_145_26), .A2 (n_0_145_32), .A3 (n_0_145_29));
NOR2_X1 i_0_145_32 (.ZN (n_0_145_32), .A1 (n_0_145_0), .A2 (n_0_145_18));
INV_X1 i_0_145_31 (.ZN (n_0_145_31), .A (n_0_145_18));
INV_X1 i_0_145_30 (.ZN (n_0_145_30), .A (n_0_145_0));
NOR2_X1 i_0_145_29 (.ZN (n_0_145_29), .A1 (n_0_145_5), .A2 (n_0_145_14));
INV_X1 i_0_145_28 (.ZN (n_0_145_28), .A (n_0_145_14));
INV_X1 i_0_145_27 (.ZN (n_0_145_27), .A (n_0_145_5));
INV_X1 i_0_145_26 (.ZN (n_0_145_26), .A (n_0_145_25));
NAND2_X1 i_0_145_25 (.ZN (n_0_145_25), .A1 (n_0_145_10), .A2 (data[6]));
NAND2_X1 i_0_145_24 (.ZN (n_0_145_24), .A1 (n_0_145_30), .A2 (n_0_145_27));
NAND3_X1 i_0_145_23 (.ZN (n_0_145_23), .A1 (n_0_145_31), .A2 (n_0_145_28), .A3 (n_0_145_10));
INV_X1 i_0_145_22 (.ZN (n_0_145_22), .A (sps__n36));
INV_X1 i_0_145_21 (.ZN (n_0_145_21), .A (sps__n7));
INV_X1 i_0_145_20 (.ZN (n_0_145_20), .A (sps__n13));
INV_X1 i_0_145_19 (.ZN (n_0_145_19), .A (address[11]));
NAND4_X1 i_0_145_18 (.ZN (n_0_145_18), .A1 (n_0_145_22), .A2 (n_0_145_21), .A3 (n_0_145_20), .A4 (n_0_145_19));
INV_X1 i_0_145_17 (.ZN (n_0_145_17), .A (sps__n61));
INV_X1 i_0_145_12 (.ZN (n_0_145_16), .A (read_signal));
INV_X1 i_0_145_11 (.ZN (n_0_145_15), .A (address[15]));
NAND4_X1 i_0_145_6 (.ZN (n_0_145_14), .A1 (n_0_145_17), .A2 (n_0_145_16), .A3 (n_0_145_15), .A4 (write_signal));
INV_X1 i_0_145_5 (.ZN (n_0_145_13), .A (sps__n113));
INV_X1 i_0_145_4 (.ZN (n_0_145_12), .A (sps__n97));
NAND3_X1 i_0_145_1 (.ZN (n_0_145_11), .A1 (n_0_145_13), .A2 (n_0_145_12), .A3 (address[2]));
INV_X1 i_0_145_0 (.ZN (n_0_145_10), .A (n_0_145_11));
INV_X1 i_0_145_16 (.ZN (n_0_145_9), .A (sps__n69));
INV_X1 i_0_145_15 (.ZN (n_0_145_8), .A (sps__n20));
INV_X1 i_0_145_14 (.ZN (n_0_145_7), .A (sps__n79));
INV_X1 i_0_145_13 (.ZN (n_0_145_6), .A (sps__n106));
NAND4_X1 i_0_145_3 (.ZN (n_0_145_5), .A1 (n_0_145_9), .A2 (n_0_145_8), .A3 (n_0_145_7), .A4 (n_0_145_6));
INV_X1 i_0_145_10 (.ZN (n_0_145_4), .A (sps__n56));
INV_X1 i_0_145_9 (.ZN (n_0_145_3), .A (sps__n27));
INV_X1 i_0_145_8 (.ZN (n_0_145_2), .A (sps__n41));
INV_X1 i_0_145_7 (.ZN (n_0_145_1), .A (sps__n93));
NAND4_X1 i_0_145_2 (.ZN (n_0_145_0), .A1 (n_0_145_4), .A2 (n_0_145_3), .A3 (n_0_145_2), .A4 (n_0_145_1));
NAND3_X1 i_0_128_31 (.ZN (n_0_128_30), .A1 (n_0_128_27), .A2 (n_0_128_28), .A3 (n_0_128_29));
NOR2_X1 i_0_128_30 (.ZN (n_0_128_29), .A1 (n_0_128_13), .A2 (n_0_128_23));
NOR2_X1 i_0_128_29 (.ZN (n_0_128_28), .A1 (n_0_128_22), .A2 (n_0_128_21));
NOR2_X1 i_0_128_28 (.ZN (n_0_128_27), .A1 (n_0_128_17), .A2 (n_0_128_20));
NOR2_X1 i_0_128_27 (.ZN (n_0_128_26), .A1 (n_0_128_17), .A2 (n_0_128_13));
NOR2_X1 i_0_128_26 (.ZN (n_0_128_25), .A1 (n_0_128_20), .A2 (n_0_128_21));
NOR2_X1 i_0_128_25 (.ZN (n_0_128_24), .A1 (n_0_128_22), .A2 (n_0_128_23));
NAND3_X1 i_0_128_24 (.ZN (n_0_128_23), .A1 (n_0_128_4), .A2 (n_0_128_2), .A3 (n_0_128_6));
NAND3_X1 i_0_128_23 (.ZN (n_0_128_22), .A1 (n_0_128_1), .A2 (n_0_128_3), .A3 (n_0_128_5));
NAND3_X1 i_0_128_22 (.ZN (n_0_128_21), .A1 (n_0_128_10), .A2 (n_0_128_8), .A3 (n_0_128_12));
NAND3_X1 i_0_128_21 (.ZN (n_0_128_20), .A1 (n_0_128_7), .A2 (n_0_128_9), .A3 (n_0_128_11));
NAND2_X1 i_0_128_20 (.ZN (n_0_128_19), .A1 (n_0_128_30), .A2 (\mem[5][6] ));
INV_X1 i_0_128_19 (.ZN (n_0_128_18), .A (sps__n114));
NAND4_X1 i_0_128_18 (.ZN (n_0_128_17), .A1 (n_0_128_18), .A2 (sps__n1), .A3 (address[2]), .A4 (sps__n97));
INV_X1 i_0_128_17 (.ZN (n_0_128_16), .A (sps__n20));
INV_X1 i_0_128_16 (.ZN (n_0_128_15), .A (sps__n79));
INV_X1 i_0_128_15 (.ZN (n_0_128_14), .A (sps__n106));
NAND3_X1 i_0_128_14 (.ZN (n_0_128_13), .A1 (n_0_128_16), .A2 (n_0_128_15), .A3 (n_0_128_14));
INV_X1 i_0_128_13 (.ZN (n_0_128_12), .A (RST));
INV_X1 i_0_128_12 (.ZN (n_0_128_11), .A (read_signal));
INV_X1 i_0_128_11 (.ZN (n_0_128_10), .A (sps__n7));
INV_X1 i_0_128_10 (.ZN (n_0_128_9), .A (sps__n13));
INV_X1 i_0_128_9 (.ZN (n_0_128_8), .A (address[15]));
INV_X1 i_0_128_8 (.ZN (n_0_128_7), .A (sps__n36));
INV_X1 i_0_128_7 (.ZN (n_0_128_6), .A (sps__n93));
INV_X1 i_0_128_6 (.ZN (n_0_128_5), .A (sps__n69));
INV_X1 i_0_128_5 (.ZN (n_0_128_4), .A (sps__n26));
INV_X1 i_0_128_4 (.ZN (n_0_128_3), .A (address[8]));
INV_X1 i_0_128_3 (.ZN (n_0_128_2), .A (address[11]));
INV_X1 i_0_128_2 (.ZN (n_0_128_1), .A (sps__n56));
NAND4_X1 i_0_128_1 (.ZN (n_0_128_0), .A1 (n_0_128_26), .A2 (n_0_128_25), .A3 (n_0_128_24), .A4 (data[6]));
NAND2_X1 i_0_128_0 (.ZN (n_0_139), .A1 (n_0_128_19), .A2 (n_0_128_0));
NAND3_X1 i_0_111_31 (.ZN (n_0_111_30), .A1 (n_0_111_27), .A2 (n_0_111_28), .A3 (n_0_111_29));
NOR2_X1 i_0_111_30 (.ZN (n_0_111_29), .A1 (n_0_111_13), .A2 (n_0_111_23));
NOR2_X1 i_0_111_29 (.ZN (n_0_111_28), .A1 (n_0_111_22), .A2 (n_0_111_21));
NOR2_X1 i_0_111_28 (.ZN (n_0_111_27), .A1 (n_0_111_17), .A2 (n_0_111_20));
NOR2_X1 i_0_111_27 (.ZN (n_0_111_26), .A1 (n_0_111_17), .A2 (n_0_111_13));
NOR2_X1 i_0_111_26 (.ZN (n_0_111_25), .A1 (n_0_111_20), .A2 (n_0_111_21));
NOR2_X1 i_0_111_25 (.ZN (n_0_111_24), .A1 (n_0_111_22), .A2 (n_0_111_23));
NAND3_X1 i_0_111_24 (.ZN (n_0_111_23), .A1 (n_0_111_4), .A2 (n_0_111_2), .A3 (n_0_111_6));
NAND3_X1 i_0_111_23 (.ZN (n_0_111_22), .A1 (n_0_111_1), .A2 (n_0_111_3), .A3 (n_0_111_5));
NAND3_X1 i_0_111_22 (.ZN (n_0_111_21), .A1 (n_0_111_10), .A2 (n_0_111_8), .A3 (n_0_111_12));
NAND3_X1 i_0_111_21 (.ZN (n_0_111_20), .A1 (n_0_111_7), .A2 (n_0_111_9), .A3 (n_0_111_11));
NAND2_X1 i_0_111_20 (.ZN (n_0_111_19), .A1 (n_0_111_30), .A2 (\mem[6][6] ));
INV_X1 i_0_111_19 (.ZN (n_0_111_18), .A (sps__n97));
NAND4_X1 i_0_111_18 (.ZN (n_0_111_17), .A1 (n_0_111_18), .A2 (sps__n1), .A3 (address[2]), .A4 (sps__n113));
INV_X1 i_0_111_17 (.ZN (n_0_111_16), .A (sps__n20));
INV_X1 i_0_111_16 (.ZN (n_0_111_15), .A (sps__n79));
INV_X1 i_0_111_15 (.ZN (n_0_111_14), .A (sps__n103));
NAND3_X1 i_0_111_14 (.ZN (n_0_111_13), .A1 (n_0_111_16), .A2 (n_0_111_15), .A3 (n_0_111_14));
INV_X1 i_0_111_13 (.ZN (n_0_111_12), .A (sps__n61));
INV_X1 i_0_111_12 (.ZN (n_0_111_11), .A (sps__n73));
INV_X1 i_0_111_11 (.ZN (n_0_111_10), .A (sps__n7));
INV_X1 i_0_111_10 (.ZN (n_0_111_9), .A (address[12]));
INV_X1 i_0_111_9 (.ZN (n_0_111_8), .A (sps__n85));
INV_X1 i_0_111_8 (.ZN (n_0_111_7), .A (sps__n36));
INV_X1 i_0_111_7 (.ZN (n_0_111_6), .A (sps__n93));
INV_X1 i_0_111_6 (.ZN (n_0_111_5), .A (sps__n69));
INV_X1 i_0_111_5 (.ZN (n_0_111_4), .A (sps__n27));
INV_X1 i_0_111_4 (.ZN (n_0_111_3), .A (sps__n41));
INV_X1 i_0_111_3 (.ZN (n_0_111_2), .A (sps__n49));
INV_X1 i_0_111_2 (.ZN (n_0_111_1), .A (sps__n56));
NAND4_X1 i_0_111_1 (.ZN (n_0_111_0), .A1 (n_0_111_26), .A2 (n_0_111_25), .A3 (n_0_111_24), .A4 (data[6]));
NAND2_X1 i_0_111_0 (.ZN (n_0_138), .A1 (n_0_111_19), .A2 (n_0_111_0));
NAND3_X1 i_0_94_27 (.ZN (n_0_94_26), .A1 (n_0_94_23), .A2 (n_0_94_24), .A3 (n_0_94_25));
NOR2_X1 i_0_94_26 (.ZN (n_0_94_25), .A1 (n_0_94_17), .A2 (n_0_94_13));
NOR2_X1 i_0_94_25 (.ZN (n_0_94_24), .A1 (n_0_94_19), .A2 (n_0_94_20));
NOR2_X1 i_0_94_24 (.ZN (n_0_94_23), .A1 (n_0_94_21), .A2 (n_0_94_22));
NAND3_X1 i_0_94_23 (.ZN (n_0_94_22), .A1 (n_0_94_4), .A2 (n_0_94_2), .A3 (n_0_94_6));
NAND3_X1 i_0_94_22 (.ZN (n_0_94_21), .A1 (n_0_94_1), .A2 (n_0_94_3), .A3 (n_0_94_5));
NAND3_X1 i_0_94_21 (.ZN (n_0_94_20), .A1 (n_0_94_10), .A2 (n_0_94_8), .A3 (n_0_94_12));
NAND3_X1 i_0_94_20 (.ZN (n_0_94_19), .A1 (n_0_94_7), .A2 (n_0_94_9), .A3 (n_0_94_11));
NAND2_X1 i_0_94_19 (.ZN (n_0_94_18), .A1 (n_0_94_26), .A2 (\mem[7][6] ));
NAND4_X1 i_0_94_18 (.ZN (n_0_94_17), .A1 (sps__n1), .A2 (address[2]), .A3 (sps__n114), .A4 (sps__n97));
INV_X1 i_0_94_17 (.ZN (n_0_94_16), .A (sps__n20));
INV_X1 i_0_94_16 (.ZN (n_0_94_15), .A (sps__n79));
INV_X1 i_0_94_15 (.ZN (n_0_94_14), .A (address[3]));
NAND3_X1 i_0_94_14 (.ZN (n_0_94_13), .A1 (n_0_94_16), .A2 (n_0_94_15), .A3 (n_0_94_14));
INV_X1 i_0_94_13 (.ZN (n_0_94_12), .A (RST));
INV_X1 i_0_94_12 (.ZN (n_0_94_11), .A (read_signal));
INV_X1 i_0_94_11 (.ZN (n_0_94_10), .A (sps__n7));
INV_X1 i_0_94_10 (.ZN (n_0_94_9), .A (sps__n13));
INV_X1 i_0_94_9 (.ZN (n_0_94_8), .A (address[15]));
INV_X1 i_0_94_8 (.ZN (n_0_94_7), .A (sps__n36));
INV_X1 i_0_94_7 (.ZN (n_0_94_6), .A (sps__n93));
INV_X1 i_0_94_6 (.ZN (n_0_94_5), .A (sps__n69));
INV_X1 i_0_94_5 (.ZN (n_0_94_4), .A (sps__n26));
INV_X1 i_0_94_4 (.ZN (n_0_94_3), .A (address[8]));
INV_X1 i_0_94_3 (.ZN (n_0_94_2), .A (address[11]));
INV_X1 i_0_94_2 (.ZN (n_0_94_1), .A (sps__n56));
NAND4_X1 i_0_94_1 (.ZN (n_0_94_0), .A1 (n_0_94_25), .A2 (n_0_94_24), .A3 (n_0_94_23), .A4 (data[6]));
NAND2_X1 i_0_94_0 (.ZN (n_0_137), .A1 (n_0_94_18), .A2 (n_0_94_0));
NAND3_X1 i_0_77_35 (.ZN (n_0_136), .A1 (n_0_77_32), .A2 (n_0_77_33), .A3 (n_0_77_34));
NAND2_X1 i_0_77_34 (.ZN (n_0_77_34), .A1 (n_0_77_23), .A2 (\mem[8][6] ));
NAND3_X1 i_0_77_29 (.ZN (n_0_77_33), .A1 (n_0_77_26), .A2 (n_0_77_31), .A3 (n_0_77_28));
NAND2_X1 i_0_77_28 (.ZN (n_0_77_32), .A1 (n_0_77_27), .A2 (\mem[8][6] ));
NOR2_X1 i_0_77_24 (.ZN (n_0_77_31), .A1 (n_0_77_18), .A2 (n_0_77_0));
INV_X1 i_0_77_23 (.ZN (n_0_77_30), .A (n_0_77_0));
INV_X1 i_0_77_22 (.ZN (n_0_77_29), .A (n_0_77_18));
INV_X1 i_0_77_21 (.ZN (n_0_77_28), .A (n_0_77_5));
NAND3_X1 i_0_77_20 (.ZN (n_0_77_27), .A1 (n_0_77_28), .A2 (n_0_77_30), .A3 (n_0_77_9));
NOR2_X1 i_0_77_19 (.ZN (n_0_77_26), .A1 (n_0_77_14), .A2 (n_0_77_24));
INV_X1 i_0_77_18 (.ZN (n_0_77_25), .A (n_0_77_14));
NAND2_X1 i_0_77_17 (.ZN (n_0_77_24), .A1 (n_0_77_9), .A2 (data[6]));
NAND2_X1 i_0_77_16 (.ZN (n_0_77_23), .A1 (n_0_77_29), .A2 (n_0_77_25));
INV_X1 i_0_77_33 (.ZN (n_0_77_22), .A (sps__n36));
INV_X1 i_0_77_32 (.ZN (n_0_77_21), .A (sps__n7));
INV_X1 i_0_77_31 (.ZN (n_0_77_20), .A (address[12]));
INV_X1 i_0_77_30 (.ZN (n_0_77_19), .A (sps__n49));
NAND4_X1 i_0_77_3 (.ZN (n_0_77_18), .A1 (n_0_77_22), .A2 (n_0_77_21), .A3 (n_0_77_20), .A4 (n_0_77_19));
INV_X1 i_0_77_27 (.ZN (n_0_77_17), .A (RST));
INV_X1 i_0_77_26 (.ZN (n_0_77_16), .A (sps__n73));
INV_X1 i_0_77_25 (.ZN (n_0_77_15), .A (sps__n85));
NAND4_X1 i_0_77_8 (.ZN (n_0_77_14), .A1 (n_0_77_17), .A2 (n_0_77_16), .A3 (n_0_77_15), .A4 (sps__n1));
INV_X1 i_0_77_15 (.ZN (n_0_77_13), .A (address[2]));
INV_X1 i_0_77_14 (.ZN (n_0_77_12), .A (sps__n114));
INV_X1 i_0_77_13 (.ZN (n_0_77_11), .A (sps__n97));
NAND3_X1 i_0_77_12 (.ZN (n_0_77_10), .A1 (n_0_77_13), .A2 (n_0_77_12), .A3 (n_0_77_11));
INV_X1 i_0_77_11 (.ZN (n_0_77_9), .A (n_0_77_10));
INV_X1 i_0_77_10 (.ZN (n_0_77_8), .A (sps__n69));
INV_X1 i_0_77_9 (.ZN (n_0_77_7), .A (sps__n20));
INV_X1 i_0_77_7 (.ZN (n_0_77_6), .A (sps__n79));
NAND4_X1 i_0_77_6 (.ZN (n_0_77_5), .A1 (n_0_77_8), .A2 (n_0_77_7), .A3 (n_0_77_6), .A4 (address[3]));
INV_X1 i_0_77_5 (.ZN (n_0_77_4), .A (sps__n56));
INV_X1 i_0_77_4 (.ZN (n_0_77_3), .A (sps__n26));
INV_X1 i_0_77_2 (.ZN (n_0_77_2), .A (address[8]));
INV_X1 i_0_77_1 (.ZN (n_0_77_1), .A (address[7]));
NAND4_X1 i_0_77_0 (.ZN (n_0_77_0), .A1 (n_0_77_4), .A2 (n_0_77_3), .A3 (n_0_77_2), .A4 (n_0_77_1));
NOR2_X1 i_0_60_34 (.ZN (n_0_60_33), .A1 (n_0_60_19), .A2 (n_0_60_0));
INV_X1 i_0_60_33 (.ZN (n_0_60_32), .A (n_0_60_0));
INV_X1 i_0_60_28 (.ZN (n_0_60_31), .A (n_0_60_19));
NAND2_X1 i_0_60_27 (.ZN (n_0_60_30), .A1 (n_0_60_29), .A2 (\mem[9][6] ));
NAND3_X1 i_0_60_23 (.ZN (n_0_60_29), .A1 (n_0_60_5), .A2 (n_0_60_32), .A3 (n_0_60_10));
NAND3_X1 i_0_60_22 (.ZN (n_0_60_28), .A1 (n_0_60_27), .A2 (n_0_60_33), .A3 (n_0_60_14));
NOR2_X1 i_0_60_21 (.ZN (n_0_60_27), .A1 (n_0_60_6), .A2 (n_0_60_26));
NAND2_X1 i_0_60_20 (.ZN (n_0_60_26), .A1 (n_0_60_10), .A2 (data[6]));
NAND2_X1 i_0_60_19 (.ZN (n_0_60_25), .A1 (n_0_60_31), .A2 (n_0_60_14));
NAND3_X1 i_0_60_18 (.ZN (n_0_135), .A1 (n_0_60_28), .A2 (n_0_60_30), .A3 (n_0_60_24));
NAND2_X1 i_0_60_17 (.ZN (n_0_60_24), .A1 (n_0_60_25), .A2 (\mem[9][6] ));
INV_X1 i_0_60_32 (.ZN (n_0_60_23), .A (sps__n36));
INV_X1 i_0_60_31 (.ZN (n_0_60_22), .A (sps__n7));
INV_X1 i_0_60_30 (.ZN (n_0_60_21), .A (address[12]));
INV_X1 i_0_60_29 (.ZN (n_0_60_20), .A (address[11]));
NAND4_X1 i_0_60_3 (.ZN (n_0_60_19), .A1 (n_0_60_23), .A2 (n_0_60_22), .A3 (n_0_60_21), .A4 (n_0_60_20));
INV_X1 i_0_60_26 (.ZN (n_0_60_18), .A (RST));
INV_X1 i_0_60_25 (.ZN (n_0_60_17), .A (sps__n73));
INV_X1 i_0_60_24 (.ZN (n_0_60_16), .A (sps__n85));
NAND4_X1 i_0_60_6 (.ZN (n_0_60_15), .A1 (n_0_60_18), .A2 (n_0_60_17), .A3 (n_0_60_16), .A4 (sps__n1));
INV_X1 i_0_60_16 (.ZN (n_0_60_14), .A (n_0_60_15));
INV_X1 i_0_60_15 (.ZN (n_0_60_13), .A (address[2]));
INV_X1 i_0_60_14 (.ZN (n_0_60_12), .A (sps__n114));
NAND3_X1 i_0_60_13 (.ZN (n_0_60_11), .A1 (n_0_60_13), .A2 (n_0_60_12), .A3 (sps__n97));
INV_X1 i_0_60_12 (.ZN (n_0_60_10), .A (n_0_60_11));
INV_X1 i_0_60_11 (.ZN (n_0_60_9), .A (sps__n69));
INV_X1 i_0_60_10 (.ZN (n_0_60_8), .A (sps__n20));
INV_X1 i_0_60_9 (.ZN (n_0_60_7), .A (sps__n79));
NAND4_X1 i_0_60_8 (.ZN (n_0_60_6), .A1 (n_0_60_9), .A2 (n_0_60_8), .A3 (n_0_60_7), .A4 (address[3]));
INV_X1 i_0_60_7 (.ZN (n_0_60_5), .A (n_0_60_6));
INV_X1 i_0_60_5 (.ZN (n_0_60_4), .A (sps__n56));
INV_X1 i_0_60_4 (.ZN (n_0_60_3), .A (sps__n26));
INV_X1 i_0_60_2 (.ZN (n_0_60_2), .A (address[8]));
INV_X1 i_0_60_1 (.ZN (n_0_60_1), .A (address[7]));
NAND4_X1 i_0_60_0 (.ZN (n_0_60_0), .A1 (n_0_60_4), .A2 (n_0_60_3), .A3 (n_0_60_2), .A4 (n_0_60_1));
NOR2_X1 i_0_43_34 (.ZN (n_0_43_33), .A1 (n_0_43_19), .A2 (n_0_43_0));
INV_X1 i_0_43_33 (.ZN (n_0_43_32), .A (n_0_43_0));
INV_X1 i_0_43_28 (.ZN (n_0_43_31), .A (n_0_43_19));
NAND2_X1 i_0_43_27 (.ZN (n_0_43_30), .A1 (n_0_43_29), .A2 (\mem[10][6] ));
NAND3_X1 i_0_43_23 (.ZN (n_0_43_29), .A1 (n_0_43_5), .A2 (n_0_43_32), .A3 (n_0_43_10));
NAND3_X1 i_0_43_22 (.ZN (n_0_43_28), .A1 (n_0_43_27), .A2 (n_0_43_33), .A3 (n_0_43_14));
NOR2_X1 i_0_43_21 (.ZN (n_0_43_27), .A1 (n_0_43_6), .A2 (n_0_43_26));
NAND2_X1 i_0_43_20 (.ZN (n_0_43_26), .A1 (n_0_43_10), .A2 (data[6]));
NAND2_X1 i_0_43_19 (.ZN (n_0_43_25), .A1 (n_0_43_31), .A2 (n_0_43_14));
NAND3_X1 i_0_43_18 (.ZN (n_0_134), .A1 (n_0_43_28), .A2 (n_0_43_30), .A3 (n_0_43_24));
NAND2_X1 i_0_43_17 (.ZN (n_0_43_24), .A1 (n_0_43_25), .A2 (\mem[10][6] ));
INV_X1 i_0_43_32 (.ZN (n_0_43_23), .A (sps__n36));
INV_X1 i_0_43_31 (.ZN (n_0_43_22), .A (sps__n7));
INV_X1 i_0_43_30 (.ZN (n_0_43_21), .A (address[12]));
INV_X1 i_0_43_29 (.ZN (n_0_43_20), .A (sps__n49));
NAND4_X1 i_0_43_3 (.ZN (n_0_43_19), .A1 (n_0_43_23), .A2 (n_0_43_22), .A3 (n_0_43_21), .A4 (n_0_43_20));
INV_X1 i_0_43_26 (.ZN (n_0_43_18), .A (sps__n61));
INV_X1 i_0_43_25 (.ZN (n_0_43_17), .A (sps__n73));
INV_X1 i_0_43_24 (.ZN (n_0_43_16), .A (sps__n85));
NAND4_X1 i_0_43_6 (.ZN (n_0_43_15), .A1 (n_0_43_18), .A2 (n_0_43_17), .A3 (n_0_43_16), .A4 (sps__n1));
INV_X1 i_0_43_16 (.ZN (n_0_43_14), .A (n_0_43_15));
INV_X1 i_0_43_15 (.ZN (n_0_43_13), .A (sps__n123));
INV_X1 i_0_43_14 (.ZN (n_0_43_12), .A (sps__n97));
NAND3_X1 i_0_43_13 (.ZN (n_0_43_11), .A1 (n_0_43_13), .A2 (n_0_43_12), .A3 (sps__n114));
INV_X1 i_0_43_12 (.ZN (n_0_43_10), .A (n_0_43_11));
INV_X1 i_0_43_11 (.ZN (n_0_43_9), .A (sps__n69));
INV_X1 i_0_43_10 (.ZN (n_0_43_8), .A (sps__n20));
INV_X1 i_0_43_9 (.ZN (n_0_43_7), .A (sps__n79));
NAND4_X1 i_0_43_8 (.ZN (n_0_43_6), .A1 (n_0_43_9), .A2 (n_0_43_8), .A3 (n_0_43_7), .A4 (sps__n103));
INV_X1 i_0_43_7 (.ZN (n_0_43_5), .A (n_0_43_6));
INV_X1 i_0_43_5 (.ZN (n_0_43_4), .A (sps__n56));
INV_X1 i_0_43_4 (.ZN (n_0_43_3), .A (sps__n27));
INV_X1 i_0_43_2 (.ZN (n_0_43_2), .A (address[8]));
INV_X1 i_0_43_1 (.ZN (n_0_43_1), .A (address[7]));
NAND4_X1 i_0_43_0 (.ZN (n_0_43_0), .A1 (n_0_43_4), .A2 (n_0_43_3), .A3 (n_0_43_2), .A4 (n_0_43_1));
NAND3_X1 i_0_26_37 (.ZN (n_0_133), .A1 (n_0_26_34), .A2 (n_0_26_35), .A3 (n_0_26_36));
NAND2_X1 i_0_26_36 (.ZN (n_0_26_36), .A1 (n_0_26_25), .A2 (\mem[0][7] ));
NAND3_X1 i_0_26_35 (.ZN (n_0_26_35), .A1 (n_0_26_27), .A2 (n_0_26_33), .A3 (n_0_26_30));
NAND2_X1 i_0_26_34 (.ZN (n_0_26_34), .A1 (n_0_26_24), .A2 (\mem[0][7] ));
NOR2_X1 i_0_26_33 (.ZN (n_0_26_33), .A1 (n_0_26_0), .A2 (n_0_26_19));
INV_X1 i_0_26_32 (.ZN (n_0_26_32), .A (n_0_26_19));
INV_X1 i_0_26_31 (.ZN (n_0_26_31), .A (n_0_26_0));
NOR2_X1 i_0_26_30 (.ZN (n_0_26_30), .A1 (n_0_26_5), .A2 (n_0_26_15));
INV_X1 i_0_26_29 (.ZN (n_0_26_29), .A (n_0_26_15));
INV_X1 i_0_26_28 (.ZN (n_0_26_28), .A (n_0_26_5));
INV_X1 i_0_26_27 (.ZN (n_0_26_27), .A (n_0_26_26));
NAND2_X1 i_0_26_26 (.ZN (n_0_26_26), .A1 (n_0_26_10), .A2 (data[7]));
NAND2_X1 i_0_26_25 (.ZN (n_0_26_25), .A1 (n_0_26_31), .A2 (n_0_26_28));
NAND3_X1 i_0_26_24 (.ZN (n_0_26_24), .A1 (n_0_26_32), .A2 (n_0_26_29), .A3 (n_0_26_10));
INV_X1 i_0_26_23 (.ZN (n_0_26_23), .A (sps__n34));
INV_X1 i_0_26_22 (.ZN (n_0_26_22), .A (sps__n9));
INV_X1 i_0_26_21 (.ZN (n_0_26_21), .A (sps__n15));
INV_X1 i_0_26_20 (.ZN (n_0_26_20), .A (sps__n51));
NAND4_X1 i_0_26_19 (.ZN (n_0_26_19), .A1 (n_0_26_23), .A2 (n_0_26_22), .A3 (n_0_26_21), .A4 (n_0_26_20));
INV_X1 i_0_26_18 (.ZN (n_0_26_18), .A (sps__n62));
INV_X1 i_0_26_17 (.ZN (n_0_26_17), .A (sps__n75));
INV_X1 i_0_26_12 (.ZN (n_0_26_16), .A (sps__n86));
NAND4_X1 i_0_26_11 (.ZN (n_0_26_15), .A1 (n_0_26_18), .A2 (n_0_26_17), .A3 (n_0_26_16), .A4 (sps__n3));
INV_X1 i_0_26_6 (.ZN (n_0_26_14), .A (sps__n122));
INV_X1 i_0_26_5 (.ZN (n_0_26_13), .A (sps__n112));
INV_X1 i_0_26_4 (.ZN (n_0_26_12), .A (sps__n99));
NAND3_X1 i_0_26_1 (.ZN (n_0_26_11), .A1 (n_0_26_14), .A2 (n_0_26_13), .A3 (n_0_26_12));
INV_X1 i_0_26_0 (.ZN (n_0_26_10), .A (n_0_26_11));
INV_X1 i_0_26_16 (.ZN (n_0_26_9), .A (address[6]));
INV_X1 i_0_26_15 (.ZN (n_0_26_8), .A (sps__n19));
INV_X1 i_0_26_14 (.ZN (n_0_26_7), .A (sps__n81));
INV_X1 i_0_26_13 (.ZN (n_0_26_6), .A (sps__n105));
NAND4_X1 i_0_26_3 (.ZN (n_0_26_5), .A1 (n_0_26_9), .A2 (n_0_26_8), .A3 (n_0_26_7), .A4 (n_0_26_6));
INV_X1 i_0_26_10 (.ZN (n_0_26_4), .A (address[10]));
INV_X1 i_0_26_9 (.ZN (n_0_26_3), .A (sps__n25));
INV_X1 i_0_26_8 (.ZN (n_0_26_2), .A (sps__n42));
INV_X1 i_0_26_7 (.ZN (n_0_26_1), .A (sps__n92));
NAND4_X1 i_0_26_2 (.ZN (n_0_26_0), .A1 (n_0_26_4), .A2 (n_0_26_3), .A3 (n_0_26_2), .A4 (n_0_26_1));
NAND3_X1 i_0_84_36 (.ZN (n_0_132), .A1 (n_0_84_33), .A2 (n_0_84_34), .A3 (n_0_84_35));
NAND2_X1 i_0_84_35 (.ZN (n_0_84_35), .A1 (n_0_84_24), .A2 (\mem[1][7] ));
NAND2_X1 i_0_84_34 (.ZN (n_0_84_34), .A1 (n_0_84_23), .A2 (\mem[1][7] ));
NAND3_X1 i_0_84_33 (.ZN (n_0_84_33), .A1 (n_0_84_26), .A2 (n_0_84_32), .A3 (n_0_84_29));
NOR2_X1 i_0_84_32 (.ZN (n_0_84_32), .A1 (n_0_84_0), .A2 (n_0_84_18));
INV_X1 i_0_84_31 (.ZN (n_0_84_31), .A (n_0_84_18));
INV_X1 i_0_84_30 (.ZN (n_0_84_30), .A (n_0_84_0));
NOR2_X1 i_0_84_29 (.ZN (n_0_84_29), .A1 (n_0_84_5), .A2 (n_0_84_14));
INV_X1 i_0_84_28 (.ZN (n_0_84_28), .A (n_0_84_14));
INV_X1 i_0_84_27 (.ZN (n_0_84_27), .A (n_0_84_5));
INV_X1 i_0_84_26 (.ZN (n_0_84_26), .A (n_0_84_25));
NAND2_X1 i_0_84_25 (.ZN (n_0_84_25), .A1 (n_0_84_10), .A2 (data[7]));
NAND2_X1 i_0_84_24 (.ZN (n_0_84_24), .A1 (n_0_84_30), .A2 (n_0_84_27));
NAND3_X1 i_0_84_23 (.ZN (n_0_84_23), .A1 (n_0_84_31), .A2 (n_0_84_28), .A3 (n_0_84_10));
INV_X1 i_0_84_22 (.ZN (n_0_84_22), .A (sps__n34));
INV_X1 i_0_84_21 (.ZN (n_0_84_21), .A (sps__n9));
INV_X1 i_0_84_20 (.ZN (n_0_84_20), .A (sps__n15));
INV_X1 i_0_84_19 (.ZN (n_0_84_19), .A (sps__n51));
NAND4_X1 i_0_84_18 (.ZN (n_0_84_18), .A1 (n_0_84_22), .A2 (n_0_84_21), .A3 (n_0_84_20), .A4 (n_0_84_19));
INV_X1 i_0_84_17 (.ZN (n_0_84_17), .A (sps__n62));
INV_X1 i_0_84_12 (.ZN (n_0_84_16), .A (sps__n75));
INV_X1 i_0_84_11 (.ZN (n_0_84_15), .A (sps__n86));
NAND4_X1 i_0_84_6 (.ZN (n_0_84_14), .A1 (n_0_84_17), .A2 (n_0_84_16), .A3 (n_0_84_15), .A4 (sps__n3));
INV_X1 i_0_84_5 (.ZN (n_0_84_13), .A (sps__n122));
INV_X1 i_0_84_4 (.ZN (n_0_84_12), .A (sps__n112));
NAND3_X1 i_0_84_1 (.ZN (n_0_84_11), .A1 (n_0_84_13), .A2 (n_0_84_12), .A3 (sps__n99));
INV_X1 i_0_84_0 (.ZN (n_0_84_10), .A (n_0_84_11));
INV_X1 i_0_84_16 (.ZN (n_0_84_9), .A (sps__n67));
INV_X1 i_0_84_15 (.ZN (n_0_84_8), .A (sps__n19));
INV_X1 i_0_84_14 (.ZN (n_0_84_7), .A (sps__n81));
INV_X1 i_0_84_13 (.ZN (n_0_84_6), .A (sps__n105));
NAND4_X1 i_0_84_3 (.ZN (n_0_84_5), .A1 (n_0_84_9), .A2 (n_0_84_8), .A3 (n_0_84_7), .A4 (n_0_84_6));
INV_X1 i_0_84_10 (.ZN (n_0_84_4), .A (sps__n55));
INV_X1 i_0_84_9 (.ZN (n_0_84_3), .A (sps__n25));
INV_X1 i_0_84_8 (.ZN (n_0_84_2), .A (sps__n42));
INV_X1 i_0_84_7 (.ZN (n_0_84_1), .A (sps__n92));
NAND4_X1 i_0_84_2 (.ZN (n_0_84_0), .A1 (n_0_84_4), .A2 (n_0_84_3), .A3 (n_0_84_2), .A4 (n_0_84_1));
NAND3_X1 i_0_178_36 (.ZN (n_0_131), .A1 (n_0_178_33), .A2 (n_0_178_34), .A3 (n_0_178_35));
NAND2_X1 i_0_178_35 (.ZN (n_0_178_35), .A1 (n_0_178_24), .A2 (\mem[2][7] ));
NAND2_X1 i_0_178_34 (.ZN (n_0_178_34), .A1 (n_0_178_23), .A2 (\mem[2][7] ));
NAND3_X1 i_0_178_33 (.ZN (n_0_178_33), .A1 (n_0_178_26), .A2 (n_0_178_32), .A3 (n_0_178_29));
NOR2_X1 i_0_178_32 (.ZN (n_0_178_32), .A1 (n_0_178_0), .A2 (n_0_178_18));
INV_X1 i_0_178_31 (.ZN (n_0_178_31), .A (n_0_178_18));
INV_X1 i_0_178_30 (.ZN (n_0_178_30), .A (n_0_178_0));
NOR2_X1 i_0_178_29 (.ZN (n_0_178_29), .A1 (n_0_178_5), .A2 (n_0_178_14));
INV_X1 i_0_178_28 (.ZN (n_0_178_28), .A (n_0_178_14));
INV_X1 i_0_178_27 (.ZN (n_0_178_27), .A (n_0_178_5));
INV_X1 i_0_178_26 (.ZN (n_0_178_26), .A (n_0_178_25));
NAND2_X1 i_0_178_25 (.ZN (n_0_178_25), .A1 (n_0_178_10), .A2 (data[7]));
NAND2_X1 i_0_178_24 (.ZN (n_0_178_24), .A1 (n_0_178_30), .A2 (n_0_178_27));
NAND3_X1 i_0_178_23 (.ZN (n_0_178_23), .A1 (n_0_178_31), .A2 (n_0_178_28), .A3 (n_0_178_10));
INV_X1 i_0_178_22 (.ZN (n_0_178_22), .A (sps__n34));
INV_X1 i_0_178_21 (.ZN (n_0_178_21), .A (sps__n9));
INV_X1 i_0_178_20 (.ZN (n_0_178_20), .A (sps__n15));
INV_X1 i_0_178_19 (.ZN (n_0_178_19), .A (sps__n51));
NAND4_X1 i_0_178_18 (.ZN (n_0_178_18), .A1 (n_0_178_22), .A2 (n_0_178_21), .A3 (n_0_178_20), .A4 (n_0_178_19));
INV_X1 i_0_178_17 (.ZN (n_0_178_17), .A (sps__n62));
INV_X1 i_0_178_12 (.ZN (n_0_178_16), .A (sps__n75));
INV_X1 i_0_178_11 (.ZN (n_0_178_15), .A (sps__n86));
NAND4_X1 i_0_178_6 (.ZN (n_0_178_14), .A1 (n_0_178_17), .A2 (n_0_178_16), .A3 (n_0_178_15), .A4 (sps__n3));
INV_X1 i_0_178_5 (.ZN (n_0_178_13), .A (sps__n122));
INV_X1 i_0_178_4 (.ZN (n_0_178_12), .A (sps__n99));
NAND3_X1 i_0_178_1 (.ZN (n_0_178_11), .A1 (n_0_178_13), .A2 (n_0_178_12), .A3 (sps__n112));
INV_X1 i_0_178_0 (.ZN (n_0_178_10), .A (n_0_178_11));
INV_X1 i_0_178_16 (.ZN (n_0_178_9), .A (address[6]));
INV_X1 i_0_178_15 (.ZN (n_0_178_8), .A (sps__n19));
INV_X1 i_0_178_14 (.ZN (n_0_178_7), .A (sps__n81));
INV_X1 i_0_178_13 (.ZN (n_0_178_6), .A (sps__n105));
NAND4_X1 i_0_178_3 (.ZN (n_0_178_5), .A1 (n_0_178_9), .A2 (n_0_178_8), .A3 (n_0_178_7), .A4 (n_0_178_6));
INV_X1 i_0_178_10 (.ZN (n_0_178_4), .A (address[10]));
INV_X1 i_0_178_9 (.ZN (n_0_178_3), .A (sps__n25));
INV_X1 i_0_178_8 (.ZN (n_0_178_2), .A (sps__n42));
INV_X1 i_0_178_7 (.ZN (n_0_178_1), .A (sps__n92));
NAND4_X1 i_0_178_2 (.ZN (n_0_178_0), .A1 (n_0_178_4), .A2 (n_0_178_3), .A3 (n_0_178_2), .A4 (n_0_178_1));
NAND3_X1 i_0_161_31 (.ZN (n_0_161_30), .A1 (n_0_161_27), .A2 (n_0_161_28), .A3 (n_0_161_29));
NOR2_X1 i_0_161_30 (.ZN (n_0_161_29), .A1 (n_0_161_13), .A2 (n_0_161_23));
NOR2_X1 i_0_161_29 (.ZN (n_0_161_28), .A1 (n_0_161_22), .A2 (n_0_161_21));
NOR2_X1 i_0_161_28 (.ZN (n_0_161_27), .A1 (n_0_161_17), .A2 (n_0_161_20));
NOR2_X1 i_0_161_27 (.ZN (n_0_161_26), .A1 (n_0_161_17), .A2 (n_0_161_13));
NOR2_X1 i_0_161_26 (.ZN (n_0_161_25), .A1 (n_0_161_20), .A2 (n_0_161_21));
NOR2_X1 i_0_161_25 (.ZN (n_0_161_24), .A1 (n_0_161_22), .A2 (n_0_161_23));
NAND3_X1 i_0_161_24 (.ZN (n_0_161_23), .A1 (n_0_161_4), .A2 (n_0_161_2), .A3 (n_0_161_6));
NAND3_X1 i_0_161_23 (.ZN (n_0_161_22), .A1 (n_0_161_1), .A2 (n_0_161_3), .A3 (n_0_161_5));
NAND3_X1 i_0_161_22 (.ZN (n_0_161_21), .A1 (n_0_161_10), .A2 (n_0_161_8), .A3 (n_0_161_12));
NAND3_X1 i_0_161_21 (.ZN (n_0_161_20), .A1 (n_0_161_7), .A2 (n_0_161_9), .A3 (n_0_161_11));
NAND2_X1 i_0_161_20 (.ZN (n_0_161_19), .A1 (n_0_161_30), .A2 (\mem[3][7] ));
INV_X1 i_0_161_19 (.ZN (n_0_161_18), .A (sps__n122));
NAND4_X1 i_0_161_18 (.ZN (n_0_161_17), .A1 (n_0_161_18), .A2 (sps__n3), .A3 (sps__n112), .A4 (sps__n99));
INV_X1 i_0_161_17 (.ZN (n_0_161_16), .A (sps__n19));
INV_X1 i_0_161_16 (.ZN (n_0_161_15), .A (sps__n81));
INV_X1 i_0_161_15 (.ZN (n_0_161_14), .A (sps__n105));
NAND3_X1 i_0_161_14 (.ZN (n_0_161_13), .A1 (n_0_161_16), .A2 (n_0_161_15), .A3 (n_0_161_14));
INV_X1 i_0_161_13 (.ZN (n_0_161_12), .A (sps__n63));
INV_X1 i_0_161_12 (.ZN (n_0_161_11), .A (sps__n75));
INV_X1 i_0_161_11 (.ZN (n_0_161_10), .A (sps__n9));
INV_X1 i_0_161_10 (.ZN (n_0_161_9), .A (sps__n15));
INV_X1 i_0_161_9 (.ZN (n_0_161_8), .A (sps__n87));
INV_X1 i_0_161_8 (.ZN (n_0_161_7), .A (sps__n34));
INV_X1 i_0_161_7 (.ZN (n_0_161_6), .A (sps__n92));
INV_X1 i_0_161_6 (.ZN (n_0_161_5), .A (address[6]));
INV_X1 i_0_161_5 (.ZN (n_0_161_4), .A (sps__n28));
INV_X1 i_0_161_4 (.ZN (n_0_161_3), .A (sps__n42));
INV_X1 i_0_161_3 (.ZN (n_0_161_2), .A (sps__n51));
INV_X1 i_0_161_2 (.ZN (n_0_161_1), .A (address[10]));
NAND4_X1 i_0_161_1 (.ZN (n_0_161_0), .A1 (n_0_161_26), .A2 (n_0_161_25), .A3 (n_0_161_24), .A4 (data[7]));
NAND2_X1 i_0_161_0 (.ZN (n_0_130), .A1 (n_0_161_19), .A2 (n_0_161_0));
NAND3_X1 i_0_144_36 (.ZN (n_0_129), .A1 (n_0_144_33), .A2 (n_0_144_34), .A3 (n_0_144_35));
NAND2_X1 i_0_144_35 (.ZN (n_0_144_35), .A1 (n_0_144_24), .A2 (\mem[4][7] ));
NAND2_X1 i_0_144_34 (.ZN (n_0_144_34), .A1 (n_0_144_23), .A2 (\mem[4][7] ));
NAND3_X1 i_0_144_33 (.ZN (n_0_144_33), .A1 (n_0_144_26), .A2 (n_0_144_32), .A3 (n_0_144_29));
NOR2_X1 i_0_144_32 (.ZN (n_0_144_32), .A1 (n_0_144_0), .A2 (n_0_144_18));
INV_X1 i_0_144_31 (.ZN (n_0_144_31), .A (n_0_144_18));
INV_X1 i_0_144_30 (.ZN (n_0_144_30), .A (n_0_144_0));
NOR2_X1 i_0_144_29 (.ZN (n_0_144_29), .A1 (n_0_144_5), .A2 (n_0_144_14));
INV_X1 i_0_144_28 (.ZN (n_0_144_28), .A (n_0_144_14));
INV_X1 i_0_144_27 (.ZN (n_0_144_27), .A (n_0_144_5));
INV_X1 i_0_144_26 (.ZN (n_0_144_26), .A (n_0_144_25));
NAND2_X1 i_0_144_25 (.ZN (n_0_144_25), .A1 (n_0_144_10), .A2 (data[7]));
NAND2_X1 i_0_144_24 (.ZN (n_0_144_24), .A1 (n_0_144_30), .A2 (n_0_144_27));
NAND3_X1 i_0_144_23 (.ZN (n_0_144_23), .A1 (n_0_144_31), .A2 (n_0_144_28), .A3 (n_0_144_10));
INV_X1 i_0_144_22 (.ZN (n_0_144_22), .A (sps__n34));
INV_X1 i_0_144_21 (.ZN (n_0_144_21), .A (sps__n9));
INV_X1 i_0_144_20 (.ZN (n_0_144_20), .A (sps__n15));
INV_X1 i_0_144_19 (.ZN (n_0_144_19), .A (sps__n50));
NAND4_X1 i_0_144_18 (.ZN (n_0_144_18), .A1 (n_0_144_22), .A2 (n_0_144_21), .A3 (n_0_144_20), .A4 (n_0_144_19));
INV_X1 i_0_144_17 (.ZN (n_0_144_17), .A (sps__n62));
INV_X1 i_0_144_12 (.ZN (n_0_144_16), .A (sps__n75));
INV_X1 i_0_144_11 (.ZN (n_0_144_15), .A (sps__n86));
NAND4_X1 i_0_144_6 (.ZN (n_0_144_14), .A1 (n_0_144_17), .A2 (n_0_144_16), .A3 (n_0_144_15), .A4 (sps__n3));
INV_X1 i_0_144_5 (.ZN (n_0_144_13), .A (sps__n112));
INV_X1 i_0_144_4 (.ZN (n_0_144_12), .A (sps__n99));
NAND3_X1 i_0_144_1 (.ZN (n_0_144_11), .A1 (n_0_144_13), .A2 (n_0_144_12), .A3 (sps__n122));
INV_X1 i_0_144_0 (.ZN (n_0_144_10), .A (n_0_144_11));
INV_X1 i_0_144_16 (.ZN (n_0_144_9), .A (address[6]));
INV_X1 i_0_144_15 (.ZN (n_0_144_8), .A (sps__n19));
INV_X1 i_0_144_14 (.ZN (n_0_144_7), .A (sps__n81));
INV_X1 i_0_144_13 (.ZN (n_0_144_6), .A (sps__n105));
NAND4_X1 i_0_144_3 (.ZN (n_0_144_5), .A1 (n_0_144_9), .A2 (n_0_144_8), .A3 (n_0_144_7), .A4 (n_0_144_6));
INV_X1 i_0_144_10 (.ZN (n_0_144_4), .A (sps__n55));
INV_X1 i_0_144_9 (.ZN (n_0_144_3), .A (sps__n28));
INV_X1 i_0_144_8 (.ZN (n_0_144_2), .A (sps__n43));
INV_X1 i_0_144_7 (.ZN (n_0_144_1), .A (sps__n92));
NAND4_X1 i_0_144_2 (.ZN (n_0_144_0), .A1 (n_0_144_4), .A2 (n_0_144_3), .A3 (n_0_144_2), .A4 (n_0_144_1));
NAND3_X1 i_0_127_31 (.ZN (n_0_127_30), .A1 (n_0_127_27), .A2 (n_0_127_28), .A3 (n_0_127_29));
NOR2_X1 i_0_127_30 (.ZN (n_0_127_29), .A1 (n_0_127_13), .A2 (n_0_127_23));
NOR2_X1 i_0_127_29 (.ZN (n_0_127_28), .A1 (n_0_127_22), .A2 (n_0_127_21));
NOR2_X1 i_0_127_28 (.ZN (n_0_127_27), .A1 (n_0_127_17), .A2 (n_0_127_20));
NOR2_X1 i_0_127_27 (.ZN (n_0_127_26), .A1 (n_0_127_17), .A2 (n_0_127_13));
NOR2_X1 i_0_127_26 (.ZN (n_0_127_25), .A1 (n_0_127_20), .A2 (n_0_127_21));
NOR2_X1 i_0_127_25 (.ZN (n_0_127_24), .A1 (n_0_127_22), .A2 (n_0_127_23));
NAND3_X1 i_0_127_24 (.ZN (n_0_127_23), .A1 (n_0_127_4), .A2 (n_0_127_2), .A3 (n_0_127_6));
NAND3_X1 i_0_127_23 (.ZN (n_0_127_22), .A1 (n_0_127_1), .A2 (n_0_127_3), .A3 (n_0_127_5));
NAND3_X1 i_0_127_22 (.ZN (n_0_127_21), .A1 (n_0_127_10), .A2 (n_0_127_8), .A3 (n_0_127_12));
NAND3_X1 i_0_127_21 (.ZN (n_0_127_20), .A1 (n_0_127_7), .A2 (n_0_127_9), .A3 (n_0_127_11));
NAND2_X1 i_0_127_20 (.ZN (n_0_127_19), .A1 (n_0_127_30), .A2 (\mem[5][7] ));
INV_X1 i_0_127_19 (.ZN (n_0_127_18), .A (sps__n112));
NAND4_X1 i_0_127_18 (.ZN (n_0_127_17), .A1 (n_0_127_18), .A2 (sps__n3), .A3 (sps__n122), .A4 (sps__n99));
INV_X1 i_0_127_17 (.ZN (n_0_127_16), .A (sps__n19));
INV_X1 i_0_127_16 (.ZN (n_0_127_15), .A (sps__n81));
INV_X1 i_0_127_15 (.ZN (n_0_127_14), .A (sps__n105));
NAND3_X1 i_0_127_14 (.ZN (n_0_127_13), .A1 (n_0_127_16), .A2 (n_0_127_15), .A3 (n_0_127_14));
INV_X1 i_0_127_13 (.ZN (n_0_127_12), .A (sps__n62));
INV_X1 i_0_127_12 (.ZN (n_0_127_11), .A (sps__n75));
INV_X1 i_0_127_11 (.ZN (n_0_127_10), .A (sps__n9));
INV_X1 i_0_127_10 (.ZN (n_0_127_9), .A (sps__n15));
INV_X1 i_0_127_9 (.ZN (n_0_127_8), .A (sps__n86));
INV_X1 i_0_127_8 (.ZN (n_0_127_7), .A (sps__n34));
INV_X1 i_0_127_7 (.ZN (n_0_127_6), .A (sps__n92));
INV_X1 i_0_127_6 (.ZN (n_0_127_5), .A (sps__n67));
INV_X1 i_0_127_5 (.ZN (n_0_127_4), .A (sps__n28));
INV_X1 i_0_127_4 (.ZN (n_0_127_3), .A (sps__n43));
INV_X1 i_0_127_3 (.ZN (n_0_127_2), .A (sps__n51));
INV_X1 i_0_127_2 (.ZN (n_0_127_1), .A (sps__n55));
NAND4_X1 i_0_127_1 (.ZN (n_0_127_0), .A1 (n_0_127_26), .A2 (n_0_127_25), .A3 (n_0_127_24), .A4 (data[7]));
NAND2_X1 i_0_127_0 (.ZN (n_0_128), .A1 (n_0_127_19), .A2 (n_0_127_0));
NAND3_X1 i_0_110_31 (.ZN (n_0_110_30), .A1 (n_0_110_27), .A2 (n_0_110_28), .A3 (n_0_110_29));
NOR2_X1 i_0_110_30 (.ZN (n_0_110_29), .A1 (n_0_110_13), .A2 (n_0_110_23));
NOR2_X1 i_0_110_29 (.ZN (n_0_110_28), .A1 (n_0_110_22), .A2 (n_0_110_21));
NOR2_X1 i_0_110_28 (.ZN (n_0_110_27), .A1 (n_0_110_17), .A2 (n_0_110_20));
NOR2_X1 i_0_110_27 (.ZN (n_0_110_26), .A1 (n_0_110_17), .A2 (n_0_110_13));
NOR2_X1 i_0_110_26 (.ZN (n_0_110_25), .A1 (n_0_110_20), .A2 (n_0_110_21));
NOR2_X1 i_0_110_25 (.ZN (n_0_110_24), .A1 (n_0_110_22), .A2 (n_0_110_23));
NAND3_X1 i_0_110_24 (.ZN (n_0_110_23), .A1 (n_0_110_4), .A2 (n_0_110_2), .A3 (n_0_110_6));
NAND3_X1 i_0_110_23 (.ZN (n_0_110_22), .A1 (n_0_110_1), .A2 (n_0_110_3), .A3 (n_0_110_5));
NAND3_X1 i_0_110_22 (.ZN (n_0_110_21), .A1 (n_0_110_10), .A2 (n_0_110_8), .A3 (n_0_110_12));
NAND3_X1 i_0_110_21 (.ZN (n_0_110_20), .A1 (n_0_110_7), .A2 (n_0_110_9), .A3 (n_0_110_11));
NAND2_X1 i_0_110_20 (.ZN (n_0_110_19), .A1 (n_0_110_30), .A2 (\mem[6][7] ));
INV_X1 i_0_110_19 (.ZN (n_0_110_18), .A (sps__n99));
NAND4_X1 i_0_110_18 (.ZN (n_0_110_17), .A1 (n_0_110_18), .A2 (sps__n3), .A3 (sps__n122), .A4 (sps__n112));
INV_X1 i_0_110_17 (.ZN (n_0_110_16), .A (sps__n19));
INV_X1 i_0_110_16 (.ZN (n_0_110_15), .A (sps__n81));
INV_X1 i_0_110_15 (.ZN (n_0_110_14), .A (sps__n105));
NAND3_X1 i_0_110_14 (.ZN (n_0_110_13), .A1 (n_0_110_16), .A2 (n_0_110_15), .A3 (n_0_110_14));
INV_X1 i_0_110_13 (.ZN (n_0_110_12), .A (sps__n62));
INV_X1 i_0_110_12 (.ZN (n_0_110_11), .A (sps__n75));
INV_X1 i_0_110_11 (.ZN (n_0_110_10), .A (sps__n9));
INV_X1 i_0_110_10 (.ZN (n_0_110_9), .A (sps__n15));
INV_X1 i_0_110_9 (.ZN (n_0_110_8), .A (sps__n86));
INV_X1 i_0_110_8 (.ZN (n_0_110_7), .A (sps__n34));
INV_X1 i_0_110_7 (.ZN (n_0_110_6), .A (sps__n92));
INV_X1 i_0_110_6 (.ZN (n_0_110_5), .A (address[6]));
INV_X1 i_0_110_5 (.ZN (n_0_110_4), .A (sps__n28));
INV_X1 i_0_110_4 (.ZN (n_0_110_3), .A (sps__n42));
INV_X1 i_0_110_3 (.ZN (n_0_110_2), .A (sps__n51));
INV_X1 i_0_110_2 (.ZN (n_0_110_1), .A (address[10]));
NAND4_X1 i_0_110_1 (.ZN (n_0_110_0), .A1 (n_0_110_26), .A2 (n_0_110_25), .A3 (n_0_110_24), .A4 (data[7]));
NAND2_X1 i_0_110_0 (.ZN (n_0_127), .A1 (n_0_110_19), .A2 (n_0_110_0));
NAND3_X1 i_0_93_27 (.ZN (n_0_93_26), .A1 (n_0_93_23), .A2 (n_0_93_24), .A3 (n_0_93_25));
NOR2_X1 i_0_93_26 (.ZN (n_0_93_25), .A1 (n_0_93_17), .A2 (n_0_93_13));
NOR2_X1 i_0_93_25 (.ZN (n_0_93_24), .A1 (n_0_93_19), .A2 (n_0_93_20));
NOR2_X1 i_0_93_24 (.ZN (n_0_93_23), .A1 (n_0_93_21), .A2 (n_0_93_22));
NAND3_X1 i_0_93_23 (.ZN (n_0_93_22), .A1 (n_0_93_4), .A2 (n_0_93_2), .A3 (n_0_93_6));
NAND3_X1 i_0_93_22 (.ZN (n_0_93_21), .A1 (n_0_93_1), .A2 (n_0_93_3), .A3 (n_0_93_5));
NAND3_X1 i_0_93_21 (.ZN (n_0_93_20), .A1 (n_0_93_10), .A2 (n_0_93_8), .A3 (n_0_93_12));
NAND3_X1 i_0_93_20 (.ZN (n_0_93_19), .A1 (n_0_93_7), .A2 (n_0_93_9), .A3 (n_0_93_11));
NAND2_X1 i_0_93_19 (.ZN (n_0_93_18), .A1 (n_0_93_26), .A2 (\mem[7][7] ));
NAND4_X1 i_0_93_18 (.ZN (n_0_93_17), .A1 (sps__n3), .A2 (sps__n122), .A3 (sps__n112), .A4 (sps__n99));
INV_X1 i_0_93_17 (.ZN (n_0_93_16), .A (sps__n19));
INV_X1 i_0_93_16 (.ZN (n_0_93_15), .A (sps__n81));
INV_X1 i_0_93_15 (.ZN (n_0_93_14), .A (sps__n105));
NAND3_X1 i_0_93_14 (.ZN (n_0_93_13), .A1 (n_0_93_16), .A2 (n_0_93_15), .A3 (n_0_93_14));
INV_X1 i_0_93_13 (.ZN (n_0_93_12), .A (sps__n62));
INV_X1 i_0_93_12 (.ZN (n_0_93_11), .A (sps__n75));
INV_X1 i_0_93_11 (.ZN (n_0_93_10), .A (sps__n9));
INV_X1 i_0_93_10 (.ZN (n_0_93_9), .A (sps__n15));
INV_X1 i_0_93_9 (.ZN (n_0_93_8), .A (sps__n86));
INV_X1 i_0_93_8 (.ZN (n_0_93_7), .A (sps__n34));
INV_X1 i_0_93_7 (.ZN (n_0_93_6), .A (sps__n92));
INV_X1 i_0_93_6 (.ZN (n_0_93_5), .A (sps__n67));
INV_X1 i_0_93_5 (.ZN (n_0_93_4), .A (sps__n28));
INV_X1 i_0_93_4 (.ZN (n_0_93_3), .A (sps__n43));
INV_X1 i_0_93_3 (.ZN (n_0_93_2), .A (sps__n51));
INV_X1 i_0_93_2 (.ZN (n_0_93_1), .A (sps__n55));
NAND4_X1 i_0_93_1 (.ZN (n_0_93_0), .A1 (n_0_93_25), .A2 (n_0_93_24), .A3 (n_0_93_23), .A4 (data[7]));
NAND2_X1 i_0_93_0 (.ZN (n_0_126), .A1 (n_0_93_18), .A2 (n_0_93_0));
NAND3_X1 i_0_76_35 (.ZN (n_0_125), .A1 (n_0_76_32), .A2 (n_0_76_33), .A3 (n_0_76_34));
NAND2_X1 i_0_76_34 (.ZN (n_0_76_34), .A1 (n_0_76_23), .A2 (\mem[8][7] ));
NAND3_X1 i_0_76_29 (.ZN (n_0_76_33), .A1 (n_0_76_26), .A2 (n_0_76_31), .A3 (n_0_76_28));
NAND2_X1 i_0_76_28 (.ZN (n_0_76_32), .A1 (n_0_76_27), .A2 (\mem[8][7] ));
NOR2_X1 i_0_76_24 (.ZN (n_0_76_31), .A1 (n_0_76_18), .A2 (n_0_76_0));
INV_X1 i_0_76_23 (.ZN (n_0_76_30), .A (n_0_76_0));
INV_X1 i_0_76_22 (.ZN (n_0_76_29), .A (n_0_76_18));
INV_X1 i_0_76_21 (.ZN (n_0_76_28), .A (n_0_76_5));
NAND3_X1 i_0_76_20 (.ZN (n_0_76_27), .A1 (n_0_76_28), .A2 (n_0_76_30), .A3 (n_0_76_9));
NOR2_X1 i_0_76_19 (.ZN (n_0_76_26), .A1 (n_0_76_14), .A2 (n_0_76_24));
INV_X1 i_0_76_18 (.ZN (n_0_76_25), .A (n_0_76_14));
NAND2_X1 i_0_76_17 (.ZN (n_0_76_24), .A1 (n_0_76_9), .A2 (data[7]));
NAND2_X1 i_0_76_16 (.ZN (n_0_76_23), .A1 (n_0_76_29), .A2 (n_0_76_25));
INV_X1 i_0_76_33 (.ZN (n_0_76_22), .A (sps__n34));
INV_X1 i_0_76_32 (.ZN (n_0_76_21), .A (sps__n9));
INV_X1 i_0_76_31 (.ZN (n_0_76_20), .A (sps__n15));
INV_X1 i_0_76_30 (.ZN (n_0_76_19), .A (sps__n51));
NAND4_X1 i_0_76_3 (.ZN (n_0_76_18), .A1 (n_0_76_22), .A2 (n_0_76_21), .A3 (n_0_76_20), .A4 (n_0_76_19));
INV_X1 i_0_76_27 (.ZN (n_0_76_17), .A (sps__n62));
INV_X1 i_0_76_26 (.ZN (n_0_76_16), .A (sps__n75));
INV_X1 i_0_76_25 (.ZN (n_0_76_15), .A (sps__n86));
NAND4_X1 i_0_76_8 (.ZN (n_0_76_14), .A1 (n_0_76_17), .A2 (n_0_76_16), .A3 (n_0_76_15), .A4 (sps__n3));
INV_X1 i_0_76_15 (.ZN (n_0_76_13), .A (sps__n122));
INV_X1 i_0_76_14 (.ZN (n_0_76_12), .A (sps__n112));
INV_X1 i_0_76_13 (.ZN (n_0_76_11), .A (sps__n99));
NAND3_X1 i_0_76_12 (.ZN (n_0_76_10), .A1 (n_0_76_13), .A2 (n_0_76_12), .A3 (n_0_76_11));
INV_X1 i_0_76_11 (.ZN (n_0_76_9), .A (n_0_76_10));
INV_X1 i_0_76_10 (.ZN (n_0_76_8), .A (address[6]));
INV_X1 i_0_76_9 (.ZN (n_0_76_7), .A (sps__n19));
INV_X1 i_0_76_7 (.ZN (n_0_76_6), .A (sps__n81));
NAND4_X1 i_0_76_6 (.ZN (n_0_76_5), .A1 (n_0_76_8), .A2 (n_0_76_7), .A3 (n_0_76_6), .A4 (sps__n105));
INV_X1 i_0_76_5 (.ZN (n_0_76_4), .A (address[10]));
INV_X1 i_0_76_4 (.ZN (n_0_76_3), .A (sps__n25));
INV_X1 i_0_76_2 (.ZN (n_0_76_2), .A (sps__n42));
INV_X1 i_0_76_1 (.ZN (n_0_76_1), .A (sps__n92));
NAND4_X1 i_0_76_0 (.ZN (n_0_76_0), .A1 (n_0_76_4), .A2 (n_0_76_3), .A3 (n_0_76_2), .A4 (n_0_76_1));
NOR2_X1 i_0_59_34 (.ZN (n_0_59_33), .A1 (n_0_59_19), .A2 (n_0_59_0));
INV_X1 i_0_59_33 (.ZN (n_0_59_32), .A (n_0_59_0));
INV_X1 i_0_59_28 (.ZN (n_0_59_31), .A (n_0_59_19));
NAND2_X1 i_0_59_27 (.ZN (n_0_59_30), .A1 (n_0_59_29), .A2 (\mem[9][7] ));
NAND3_X1 i_0_59_23 (.ZN (n_0_59_29), .A1 (n_0_59_5), .A2 (n_0_59_32), .A3 (n_0_59_10));
NAND3_X1 i_0_59_22 (.ZN (n_0_59_28), .A1 (n_0_59_27), .A2 (n_0_59_33), .A3 (n_0_59_14));
NOR2_X1 i_0_59_21 (.ZN (n_0_59_27), .A1 (n_0_59_6), .A2 (n_0_59_26));
NAND2_X1 i_0_59_20 (.ZN (n_0_59_26), .A1 (n_0_59_10), .A2 (data[7]));
NAND2_X1 i_0_59_19 (.ZN (n_0_59_25), .A1 (n_0_59_31), .A2 (n_0_59_14));
NAND3_X1 i_0_59_18 (.ZN (n_0_124), .A1 (n_0_59_28), .A2 (n_0_59_30), .A3 (n_0_59_24));
NAND2_X1 i_0_59_17 (.ZN (n_0_59_24), .A1 (n_0_59_25), .A2 (\mem[9][7] ));
INV_X1 i_0_59_32 (.ZN (n_0_59_23), .A (sps__n34));
INV_X1 i_0_59_31 (.ZN (n_0_59_22), .A (sps__n9));
INV_X1 i_0_59_30 (.ZN (n_0_59_21), .A (sps__n15));
INV_X1 i_0_59_29 (.ZN (n_0_59_20), .A (sps__n51));
NAND4_X1 i_0_59_3 (.ZN (n_0_59_19), .A1 (n_0_59_23), .A2 (n_0_59_22), .A3 (n_0_59_21), .A4 (n_0_59_20));
INV_X1 i_0_59_26 (.ZN (n_0_59_18), .A (sps__n62));
INV_X1 i_0_59_25 (.ZN (n_0_59_17), .A (sps__n75));
INV_X1 i_0_59_24 (.ZN (n_0_59_16), .A (sps__n86));
NAND4_X1 i_0_59_6 (.ZN (n_0_59_15), .A1 (n_0_59_18), .A2 (n_0_59_17), .A3 (n_0_59_16), .A4 (sps__n3));
INV_X1 i_0_59_16 (.ZN (n_0_59_14), .A (n_0_59_15));
INV_X1 i_0_59_15 (.ZN (n_0_59_13), .A (sps__n122));
INV_X1 i_0_59_14 (.ZN (n_0_59_12), .A (sps__n112));
NAND3_X1 i_0_59_13 (.ZN (n_0_59_11), .A1 (n_0_59_13), .A2 (n_0_59_12), .A3 (sps__n99));
INV_X1 i_0_59_12 (.ZN (n_0_59_10), .A (n_0_59_11));
INV_X1 i_0_59_11 (.ZN (n_0_59_9), .A (address[6]));
INV_X1 i_0_59_10 (.ZN (n_0_59_8), .A (sps__n19));
INV_X1 i_0_59_9 (.ZN (n_0_59_7), .A (sps__n81));
NAND4_X1 i_0_59_8 (.ZN (n_0_59_6), .A1 (n_0_59_9), .A2 (n_0_59_8), .A3 (n_0_59_7), .A4 (sps__n105));
INV_X1 i_0_59_7 (.ZN (n_0_59_5), .A (n_0_59_6));
INV_X1 i_0_59_5 (.ZN (n_0_59_4), .A (address[10]));
INV_X1 i_0_59_4 (.ZN (n_0_59_3), .A (sps__n25));
INV_X1 i_0_59_2 (.ZN (n_0_59_2), .A (sps__n42));
INV_X1 i_0_59_1 (.ZN (n_0_59_1), .A (sps__n92));
NAND4_X1 i_0_59_0 (.ZN (n_0_59_0), .A1 (n_0_59_4), .A2 (n_0_59_3), .A3 (n_0_59_2), .A4 (n_0_59_1));
NOR2_X1 i_0_25_34 (.ZN (n_0_25_33), .A1 (n_0_25_19), .A2 (n_0_25_0));
INV_X1 i_0_25_33 (.ZN (n_0_25_32), .A (n_0_25_0));
INV_X1 i_0_25_28 (.ZN (n_0_25_31), .A (n_0_25_19));
NAND2_X1 i_0_25_27 (.ZN (n_0_25_30), .A1 (n_0_25_29), .A2 (\mem[10][7] ));
NAND3_X1 i_0_25_23 (.ZN (n_0_25_29), .A1 (n_0_25_5), .A2 (n_0_25_32), .A3 (n_0_25_10));
NAND3_X1 i_0_25_22 (.ZN (n_0_25_28), .A1 (n_0_25_27), .A2 (n_0_25_33), .A3 (n_0_25_14));
NOR2_X1 i_0_25_21 (.ZN (n_0_25_27), .A1 (n_0_25_6), .A2 (n_0_25_26));
NAND2_X1 i_0_25_20 (.ZN (n_0_25_26), .A1 (n_0_25_10), .A2 (data[7]));
NAND2_X1 i_0_25_19 (.ZN (n_0_25_25), .A1 (n_0_25_31), .A2 (n_0_25_14));
NAND3_X1 i_0_25_18 (.ZN (n_0_123), .A1 (n_0_25_28), .A2 (n_0_25_30), .A3 (n_0_25_24));
NAND2_X1 i_0_25_17 (.ZN (n_0_25_24), .A1 (n_0_25_25), .A2 (\mem[10][7] ));
INV_X1 i_0_25_32 (.ZN (n_0_25_23), .A (sps__n34));
INV_X1 i_0_25_31 (.ZN (n_0_25_22), .A (sps__n9));
INV_X1 i_0_25_30 (.ZN (n_0_25_21), .A (sps__n15));
INV_X1 i_0_25_29 (.ZN (n_0_25_20), .A (sps__n51));
NAND4_X1 i_0_25_3 (.ZN (n_0_25_19), .A1 (n_0_25_23), .A2 (n_0_25_22), .A3 (n_0_25_21), .A4 (n_0_25_20));
INV_X1 i_0_25_26 (.ZN (n_0_25_18), .A (sps__n62));
INV_X1 i_0_25_25 (.ZN (n_0_25_17), .A (sps__n75));
INV_X1 i_0_25_24 (.ZN (n_0_25_16), .A (sps__n86));
NAND4_X1 i_0_25_6 (.ZN (n_0_25_15), .A1 (n_0_25_18), .A2 (n_0_25_17), .A3 (n_0_25_16), .A4 (sps__n3));
INV_X1 i_0_25_16 (.ZN (n_0_25_14), .A (n_0_25_15));
INV_X1 i_0_25_15 (.ZN (n_0_25_13), .A (sps__n122));
INV_X1 i_0_25_14 (.ZN (n_0_25_12), .A (sps__n99));
NAND3_X1 i_0_25_13 (.ZN (n_0_25_11), .A1 (n_0_25_13), .A2 (n_0_25_12), .A3 (sps__n112));
INV_X1 i_0_25_12 (.ZN (n_0_25_10), .A (n_0_25_11));
INV_X1 i_0_25_11 (.ZN (n_0_25_9), .A (address[6]));
INV_X1 i_0_25_10 (.ZN (n_0_25_8), .A (sps__n19));
INV_X1 i_0_25_9 (.ZN (n_0_25_7), .A (sps__n81));
NAND4_X1 i_0_25_8 (.ZN (n_0_25_6), .A1 (n_0_25_9), .A2 (n_0_25_8), .A3 (n_0_25_7), .A4 (sps__n105));
INV_X1 i_0_25_7 (.ZN (n_0_25_5), .A (n_0_25_6));
INV_X1 i_0_25_5 (.ZN (n_0_25_4), .A (sps__n55));
INV_X1 i_0_25_4 (.ZN (n_0_25_3), .A (sps__n28));
INV_X1 i_0_25_2 (.ZN (n_0_25_2), .A (sps__n43));
INV_X1 i_0_25_1 (.ZN (n_0_25_1), .A (sps__n92));
NAND4_X1 i_0_25_0 (.ZN (n_0_25_0), .A1 (n_0_25_4), .A2 (n_0_25_3), .A3 (n_0_25_2), .A4 (n_0_25_1));
NAND3_X1 i_0_2_37 (.ZN (n_0_122), .A1 (n_0_2_34), .A2 (n_0_2_35), .A3 (n_0_2_36));
NAND2_X1 i_0_2_36 (.ZN (n_0_2_36), .A1 (n_0_2_25), .A2 (\mem[0][8] ));
NAND3_X1 i_0_2_35 (.ZN (n_0_2_35), .A1 (n_0_2_27), .A2 (n_0_2_33), .A3 (n_0_2_30));
NAND2_X1 i_0_2_34 (.ZN (n_0_2_34), .A1 (n_0_2_24), .A2 (\mem[0][8] ));
NOR2_X1 i_0_2_33 (.ZN (n_0_2_33), .A1 (n_0_2_0), .A2 (n_0_2_19));
INV_X1 i_0_2_32 (.ZN (n_0_2_32), .A (n_0_2_19));
INV_X1 i_0_2_31 (.ZN (n_0_2_31), .A (n_0_2_0));
NOR2_X1 i_0_2_30 (.ZN (n_0_2_30), .A1 (n_0_2_5), .A2 (n_0_2_15));
INV_X1 i_0_2_29 (.ZN (n_0_2_29), .A (n_0_2_15));
INV_X1 i_0_2_28 (.ZN (n_0_2_28), .A (n_0_2_5));
INV_X1 i_0_2_27 (.ZN (n_0_2_27), .A (n_0_2_26));
NAND2_X1 i_0_2_26 (.ZN (n_0_2_26), .A1 (n_0_2_10), .A2 (data[8]));
NAND2_X1 i_0_2_25 (.ZN (n_0_2_25), .A1 (n_0_2_31), .A2 (n_0_2_28));
NAND3_X1 i_0_2_24 (.ZN (n_0_2_24), .A1 (n_0_2_32), .A2 (n_0_2_29), .A3 (n_0_2_10));
INV_X1 i_0_2_23 (.ZN (n_0_2_23), .A (sps__n34));
INV_X1 i_0_2_22 (.ZN (n_0_2_22), .A (sps__n9));
INV_X1 i_0_2_21 (.ZN (n_0_2_21), .A (sps__n15));
INV_X1 i_0_2_20 (.ZN (n_0_2_20), .A (sps__n50));
NAND4_X1 i_0_2_19 (.ZN (n_0_2_19), .A1 (n_0_2_23), .A2 (n_0_2_22), .A3 (n_0_2_21), .A4 (n_0_2_20));
INV_X1 i_0_2_18 (.ZN (n_0_2_18), .A (sps__n62));
INV_X1 i_0_2_17 (.ZN (n_0_2_17), .A (sps__n75));
INV_X1 i_0_2_12 (.ZN (n_0_2_16), .A (sps__n87));
NAND4_X1 i_0_2_11 (.ZN (n_0_2_15), .A1 (n_0_2_18), .A2 (n_0_2_17), .A3 (n_0_2_16), .A4 (sps__n3));
INV_X1 i_0_2_6 (.ZN (n_0_2_14), .A (sps__n122));
INV_X1 i_0_2_5 (.ZN (n_0_2_13), .A (sps__n112));
INV_X1 i_0_2_4 (.ZN (n_0_2_12), .A (sps__n99));
NAND3_X1 i_0_2_1 (.ZN (n_0_2_11), .A1 (n_0_2_14), .A2 (n_0_2_13), .A3 (n_0_2_12));
INV_X1 i_0_2_0 (.ZN (n_0_2_10), .A (n_0_2_11));
INV_X1 i_0_2_16 (.ZN (n_0_2_9), .A (sps__n67));
INV_X1 i_0_2_15 (.ZN (n_0_2_8), .A (sps__n19));
INV_X1 i_0_2_14 (.ZN (n_0_2_7), .A (sps__n81));
INV_X1 i_0_2_13 (.ZN (n_0_2_6), .A (sps__n104));
NAND4_X1 i_0_2_3 (.ZN (n_0_2_5), .A1 (n_0_2_9), .A2 (n_0_2_8), .A3 (n_0_2_7), .A4 (n_0_2_6));
INV_X1 i_0_2_10 (.ZN (n_0_2_4), .A (sps__n55));
INV_X1 i_0_2_9 (.ZN (n_0_2_3), .A (sps__n26));
INV_X1 i_0_2_8 (.ZN (n_0_2_2), .A (sps__n43));
INV_X1 i_0_2_7 (.ZN (n_0_2_1), .A (sps__n91));
NAND4_X1 i_0_2_2 (.ZN (n_0_2_0), .A1 (n_0_2_4), .A2 (n_0_2_3), .A3 (n_0_2_2), .A4 (n_0_2_1));
NAND3_X1 i_0_135_36 (.ZN (n_0_121), .A1 (n_0_135_33), .A2 (n_0_135_34), .A3 (n_0_135_35));
NAND2_X1 i_0_135_35 (.ZN (n_0_135_35), .A1 (n_0_135_24), .A2 (\mem[1][8] ));
NAND2_X1 i_0_135_34 (.ZN (n_0_135_34), .A1 (n_0_135_23), .A2 (\mem[1][8] ));
NAND3_X1 i_0_135_33 (.ZN (n_0_135_33), .A1 (n_0_135_26), .A2 (n_0_135_32), .A3 (n_0_135_29));
NOR2_X1 i_0_135_32 (.ZN (n_0_135_32), .A1 (n_0_135_0), .A2 (n_0_135_18));
INV_X1 i_0_135_31 (.ZN (n_0_135_31), .A (n_0_135_18));
INV_X1 i_0_135_30 (.ZN (n_0_135_30), .A (n_0_135_0));
NOR2_X1 i_0_135_29 (.ZN (n_0_135_29), .A1 (n_0_135_5), .A2 (n_0_135_14));
INV_X1 i_0_135_28 (.ZN (n_0_135_28), .A (n_0_135_14));
INV_X1 i_0_135_27 (.ZN (n_0_135_27), .A (n_0_135_5));
INV_X1 i_0_135_26 (.ZN (n_0_135_26), .A (n_0_135_25));
NAND2_X1 i_0_135_25 (.ZN (n_0_135_25), .A1 (n_0_135_10), .A2 (data[8]));
NAND2_X1 i_0_135_24 (.ZN (n_0_135_24), .A1 (n_0_135_30), .A2 (n_0_135_27));
NAND3_X1 i_0_135_23 (.ZN (n_0_135_23), .A1 (n_0_135_31), .A2 (n_0_135_28), .A3 (n_0_135_10));
INV_X1 i_0_135_22 (.ZN (n_0_135_22), .A (sps__n34));
INV_X1 i_0_135_21 (.ZN (n_0_135_21), .A (sps__n8));
INV_X1 i_0_135_20 (.ZN (n_0_135_20), .A (sps__n14));
INV_X1 i_0_135_19 (.ZN (n_0_135_19), .A (sps__n50));
NAND4_X1 i_0_135_18 (.ZN (n_0_135_18), .A1 (n_0_135_22), .A2 (n_0_135_21), .A3 (n_0_135_20), .A4 (n_0_135_19));
INV_X1 i_0_135_17 (.ZN (n_0_135_17), .A (sps__n63));
INV_X1 i_0_135_12 (.ZN (n_0_135_16), .A (sps__n75));
INV_X1 i_0_135_11 (.ZN (n_0_135_15), .A (sps__n87));
NAND4_X1 i_0_135_6 (.ZN (n_0_135_14), .A1 (n_0_135_17), .A2 (n_0_135_16), .A3 (n_0_135_15), .A4 (sps__n3));
INV_X1 i_0_135_5 (.ZN (n_0_135_13), .A (sps__n122));
INV_X1 i_0_135_4 (.ZN (n_0_135_12), .A (sps__n112));
NAND3_X1 i_0_135_1 (.ZN (n_0_135_11), .A1 (n_0_135_13), .A2 (n_0_135_12), .A3 (sps__n99));
INV_X1 i_0_135_0 (.ZN (n_0_135_10), .A (n_0_135_11));
INV_X1 i_0_135_16 (.ZN (n_0_135_9), .A (sps__n67));
INV_X1 i_0_135_15 (.ZN (n_0_135_8), .A (sps__n19));
INV_X1 i_0_135_14 (.ZN (n_0_135_7), .A (sps__n81));
INV_X1 i_0_135_13 (.ZN (n_0_135_6), .A (sps__n104));
NAND4_X1 i_0_135_3 (.ZN (n_0_135_5), .A1 (n_0_135_9), .A2 (n_0_135_8), .A3 (n_0_135_7), .A4 (n_0_135_6));
INV_X1 i_0_135_10 (.ZN (n_0_135_4), .A (sps__n57));
INV_X1 i_0_135_9 (.ZN (n_0_135_3), .A (sps__n26));
INV_X1 i_0_135_8 (.ZN (n_0_135_2), .A (sps__n43));
INV_X1 i_0_135_7 (.ZN (n_0_135_1), .A (sps__n91));
NAND4_X1 i_0_135_2 (.ZN (n_0_135_0), .A1 (n_0_135_4), .A2 (n_0_135_3), .A3 (n_0_135_2), .A4 (n_0_135_1));
NAND3_X1 i_0_177_36 (.ZN (n_0_120), .A1 (n_0_177_33), .A2 (n_0_177_34), .A3 (n_0_177_35));
NAND2_X1 i_0_177_35 (.ZN (n_0_177_35), .A1 (n_0_177_24), .A2 (\mem[2][8] ));
NAND2_X1 i_0_177_34 (.ZN (n_0_177_34), .A1 (n_0_177_23), .A2 (\mem[2][8] ));
NAND3_X1 i_0_177_33 (.ZN (n_0_177_33), .A1 (n_0_177_26), .A2 (n_0_177_32), .A3 (n_0_177_29));
NOR2_X1 i_0_177_32 (.ZN (n_0_177_32), .A1 (n_0_177_0), .A2 (n_0_177_18));
INV_X1 i_0_177_31 (.ZN (n_0_177_31), .A (n_0_177_18));
INV_X1 i_0_177_30 (.ZN (n_0_177_30), .A (n_0_177_0));
NOR2_X1 i_0_177_29 (.ZN (n_0_177_29), .A1 (n_0_177_5), .A2 (n_0_177_14));
INV_X1 i_0_177_28 (.ZN (n_0_177_28), .A (n_0_177_14));
INV_X1 i_0_177_27 (.ZN (n_0_177_27), .A (n_0_177_5));
INV_X1 i_0_177_26 (.ZN (n_0_177_26), .A (n_0_177_25));
NAND2_X1 i_0_177_25 (.ZN (n_0_177_25), .A1 (n_0_177_10), .A2 (data[8]));
NAND2_X1 i_0_177_24 (.ZN (n_0_177_24), .A1 (n_0_177_30), .A2 (n_0_177_27));
NAND3_X1 i_0_177_23 (.ZN (n_0_177_23), .A1 (n_0_177_31), .A2 (n_0_177_28), .A3 (n_0_177_10));
INV_X1 i_0_177_22 (.ZN (n_0_177_22), .A (sps__n34));
INV_X1 i_0_177_21 (.ZN (n_0_177_21), .A (sps__n9));
INV_X1 i_0_177_20 (.ZN (n_0_177_20), .A (sps__n15));
INV_X1 i_0_177_19 (.ZN (n_0_177_19), .A (sps__n51));
NAND4_X1 i_0_177_18 (.ZN (n_0_177_18), .A1 (n_0_177_22), .A2 (n_0_177_21), .A3 (n_0_177_20), .A4 (n_0_177_19));
INV_X1 i_0_177_17 (.ZN (n_0_177_17), .A (sps__n62));
INV_X1 i_0_177_12 (.ZN (n_0_177_16), .A (sps__n75));
INV_X1 i_0_177_11 (.ZN (n_0_177_15), .A (sps__n86));
NAND4_X1 i_0_177_6 (.ZN (n_0_177_14), .A1 (n_0_177_17), .A2 (n_0_177_16), .A3 (n_0_177_15), .A4 (sps__n3));
INV_X1 i_0_177_5 (.ZN (n_0_177_13), .A (sps__n122));
INV_X1 i_0_177_4 (.ZN (n_0_177_12), .A (sps__n99));
NAND3_X1 i_0_177_1 (.ZN (n_0_177_11), .A1 (n_0_177_13), .A2 (n_0_177_12), .A3 (sps__n112));
INV_X1 i_0_177_0 (.ZN (n_0_177_10), .A (n_0_177_11));
INV_X1 i_0_177_16 (.ZN (n_0_177_9), .A (sps__n67));
INV_X1 i_0_177_15 (.ZN (n_0_177_8), .A (sps__n19));
INV_X1 i_0_177_14 (.ZN (n_0_177_7), .A (sps__n81));
INV_X1 i_0_177_13 (.ZN (n_0_177_6), .A (sps__n104));
NAND4_X1 i_0_177_3 (.ZN (n_0_177_5), .A1 (n_0_177_9), .A2 (n_0_177_8), .A3 (n_0_177_7), .A4 (n_0_177_6));
INV_X1 i_0_177_10 (.ZN (n_0_177_4), .A (sps__n55));
INV_X1 i_0_177_9 (.ZN (n_0_177_3), .A (sps__n28));
INV_X1 i_0_177_8 (.ZN (n_0_177_2), .A (sps__n43));
INV_X1 i_0_177_7 (.ZN (n_0_177_1), .A (sps__n92));
NAND4_X1 i_0_177_2 (.ZN (n_0_177_0), .A1 (n_0_177_4), .A2 (n_0_177_3), .A3 (n_0_177_2), .A4 (n_0_177_1));
NAND3_X1 i_0_160_31 (.ZN (n_0_160_30), .A1 (n_0_160_27), .A2 (n_0_160_28), .A3 (n_0_160_29));
NOR2_X1 i_0_160_30 (.ZN (n_0_160_29), .A1 (n_0_160_13), .A2 (n_0_160_23));
NOR2_X1 i_0_160_29 (.ZN (n_0_160_28), .A1 (n_0_160_22), .A2 (n_0_160_21));
NOR2_X1 i_0_160_28 (.ZN (n_0_160_27), .A1 (n_0_160_17), .A2 (n_0_160_20));
NOR2_X1 i_0_160_27 (.ZN (n_0_160_26), .A1 (n_0_160_17), .A2 (n_0_160_13));
NOR2_X1 i_0_160_26 (.ZN (n_0_160_25), .A1 (n_0_160_20), .A2 (n_0_160_21));
NOR2_X1 i_0_160_25 (.ZN (n_0_160_24), .A1 (n_0_160_22), .A2 (n_0_160_23));
NAND3_X1 i_0_160_24 (.ZN (n_0_160_23), .A1 (n_0_160_4), .A2 (n_0_160_2), .A3 (n_0_160_6));
NAND3_X1 i_0_160_23 (.ZN (n_0_160_22), .A1 (n_0_160_1), .A2 (n_0_160_3), .A3 (n_0_160_5));
NAND3_X1 i_0_160_22 (.ZN (n_0_160_21), .A1 (n_0_160_10), .A2 (n_0_160_8), .A3 (n_0_160_12));
NAND3_X1 i_0_160_21 (.ZN (n_0_160_20), .A1 (n_0_160_7), .A2 (n_0_160_9), .A3 (n_0_160_11));
NAND2_X1 i_0_160_20 (.ZN (n_0_160_19), .A1 (n_0_160_30), .A2 (\mem[3][8] ));
INV_X1 i_0_160_19 (.ZN (n_0_160_18), .A (sps__n122));
NAND4_X1 i_0_160_18 (.ZN (n_0_160_17), .A1 (n_0_160_18), .A2 (sps__n3), .A3 (sps__n112), .A4 (sps__n99));
INV_X1 i_0_160_17 (.ZN (n_0_160_16), .A (sps__n19));
INV_X1 i_0_160_16 (.ZN (n_0_160_15), .A (sps__n81));
INV_X1 i_0_160_15 (.ZN (n_0_160_14), .A (sps__n105));
NAND3_X1 i_0_160_14 (.ZN (n_0_160_13), .A1 (n_0_160_16), .A2 (n_0_160_15), .A3 (n_0_160_14));
INV_X1 i_0_160_13 (.ZN (n_0_160_12), .A (sps__n63));
INV_X1 i_0_160_12 (.ZN (n_0_160_11), .A (sps__n75));
INV_X1 i_0_160_11 (.ZN (n_0_160_10), .A (sps__n9));
INV_X1 i_0_160_10 (.ZN (n_0_160_9), .A (sps__n15));
INV_X1 i_0_160_9 (.ZN (n_0_160_8), .A (sps__n87));
INV_X1 i_0_160_8 (.ZN (n_0_160_7), .A (sps__n34));
INV_X1 i_0_160_7 (.ZN (n_0_160_6), .A (sps__n92));
INV_X1 i_0_160_6 (.ZN (n_0_160_5), .A (sps__n67));
INV_X1 i_0_160_5 (.ZN (n_0_160_4), .A (sps__n28));
INV_X1 i_0_160_4 (.ZN (n_0_160_3), .A (sps__n43));
INV_X1 i_0_160_3 (.ZN (n_0_160_2), .A (sps__n51));
INV_X1 i_0_160_2 (.ZN (n_0_160_1), .A (sps__n55));
NAND4_X1 i_0_160_1 (.ZN (n_0_160_0), .A1 (n_0_160_26), .A2 (n_0_160_25), .A3 (n_0_160_24), .A4 (data[8]));
NAND2_X1 i_0_160_0 (.ZN (n_0_119), .A1 (n_0_160_19), .A2 (n_0_160_0));
NAND3_X1 i_0_143_36 (.ZN (n_0_118), .A1 (n_0_143_33), .A2 (n_0_143_34), .A3 (n_0_143_35));
NAND2_X1 i_0_143_35 (.ZN (n_0_143_35), .A1 (n_0_143_24), .A2 (\mem[4][8] ));
NAND2_X1 i_0_143_34 (.ZN (n_0_143_34), .A1 (n_0_143_23), .A2 (\mem[4][8] ));
NAND3_X1 i_0_143_33 (.ZN (n_0_143_33), .A1 (n_0_143_26), .A2 (n_0_143_32), .A3 (n_0_143_29));
NOR2_X1 i_0_143_32 (.ZN (n_0_143_32), .A1 (n_0_143_0), .A2 (n_0_143_18));
INV_X1 i_0_143_31 (.ZN (n_0_143_31), .A (n_0_143_18));
INV_X1 i_0_143_30 (.ZN (n_0_143_30), .A (n_0_143_0));
NOR2_X1 i_0_143_29 (.ZN (n_0_143_29), .A1 (n_0_143_5), .A2 (n_0_143_14));
INV_X1 i_0_143_28 (.ZN (n_0_143_28), .A (n_0_143_14));
INV_X1 i_0_143_27 (.ZN (n_0_143_27), .A (n_0_143_5));
INV_X1 i_0_143_26 (.ZN (n_0_143_26), .A (n_0_143_25));
NAND2_X1 i_0_143_25 (.ZN (n_0_143_25), .A1 (n_0_143_10), .A2 (data[8]));
NAND2_X1 i_0_143_24 (.ZN (n_0_143_24), .A1 (n_0_143_30), .A2 (n_0_143_27));
NAND3_X1 i_0_143_23 (.ZN (n_0_143_23), .A1 (n_0_143_31), .A2 (n_0_143_28), .A3 (n_0_143_10));
INV_X1 i_0_143_22 (.ZN (n_0_143_22), .A (sps__n34));
INV_X1 i_0_143_21 (.ZN (n_0_143_21), .A (sps__n8));
INV_X1 i_0_143_20 (.ZN (n_0_143_20), .A (sps__n14));
INV_X1 i_0_143_19 (.ZN (n_0_143_19), .A (sps__n50));
NAND4_X1 i_0_143_18 (.ZN (n_0_143_18), .A1 (n_0_143_22), .A2 (n_0_143_21), .A3 (n_0_143_20), .A4 (n_0_143_19));
INV_X1 i_0_143_17 (.ZN (n_0_143_17), .A (sps__n63));
INV_X1 i_0_143_12 (.ZN (n_0_143_16), .A (sps__n75));
INV_X1 i_0_143_11 (.ZN (n_0_143_15), .A (sps__n87));
NAND4_X1 i_0_143_6 (.ZN (n_0_143_14), .A1 (n_0_143_17), .A2 (n_0_143_16), .A3 (n_0_143_15), .A4 (sps__n3));
INV_X1 i_0_143_5 (.ZN (n_0_143_13), .A (sps__n112));
INV_X1 i_0_143_4 (.ZN (n_0_143_12), .A (sps__n99));
NAND3_X1 i_0_143_1 (.ZN (n_0_143_11), .A1 (n_0_143_13), .A2 (n_0_143_12), .A3 (sps__n122));
INV_X1 i_0_143_0 (.ZN (n_0_143_10), .A (n_0_143_11));
INV_X1 i_0_143_16 (.ZN (n_0_143_9), .A (sps__n67));
INV_X1 i_0_143_15 (.ZN (n_0_143_8), .A (sps__n19));
INV_X1 i_0_143_14 (.ZN (n_0_143_7), .A (sps__n81));
INV_X1 i_0_143_13 (.ZN (n_0_143_6), .A (sps__n104));
NAND4_X1 i_0_143_3 (.ZN (n_0_143_5), .A1 (n_0_143_9), .A2 (n_0_143_8), .A3 (n_0_143_7), .A4 (n_0_143_6));
INV_X1 i_0_143_10 (.ZN (n_0_143_4), .A (sps__n57));
INV_X1 i_0_143_9 (.ZN (n_0_143_3), .A (sps__n26));
INV_X1 i_0_143_8 (.ZN (n_0_143_2), .A (sps__n43));
INV_X1 i_0_143_7 (.ZN (n_0_143_1), .A (sps__n91));
NAND4_X1 i_0_143_2 (.ZN (n_0_143_0), .A1 (n_0_143_4), .A2 (n_0_143_3), .A3 (n_0_143_2), .A4 (n_0_143_1));
NAND3_X1 i_0_126_31 (.ZN (n_0_126_30), .A1 (n_0_126_27), .A2 (n_0_126_28), .A3 (n_0_126_29));
NOR2_X1 i_0_126_30 (.ZN (n_0_126_29), .A1 (n_0_126_13), .A2 (n_0_126_23));
NOR2_X1 i_0_126_29 (.ZN (n_0_126_28), .A1 (n_0_126_22), .A2 (n_0_126_21));
NOR2_X1 i_0_126_28 (.ZN (n_0_126_27), .A1 (n_0_126_17), .A2 (n_0_126_20));
NOR2_X1 i_0_126_27 (.ZN (n_0_126_26), .A1 (n_0_126_17), .A2 (n_0_126_13));
NOR2_X1 i_0_126_26 (.ZN (n_0_126_25), .A1 (n_0_126_20), .A2 (n_0_126_21));
NOR2_X1 i_0_126_25 (.ZN (n_0_126_24), .A1 (n_0_126_22), .A2 (n_0_126_23));
NAND3_X1 i_0_126_24 (.ZN (n_0_126_23), .A1 (n_0_126_4), .A2 (n_0_126_2), .A3 (n_0_126_6));
NAND3_X1 i_0_126_23 (.ZN (n_0_126_22), .A1 (n_0_126_1), .A2 (n_0_126_3), .A3 (n_0_126_5));
NAND3_X1 i_0_126_22 (.ZN (n_0_126_21), .A1 (n_0_126_10), .A2 (n_0_126_8), .A3 (n_0_126_12));
NAND3_X1 i_0_126_21 (.ZN (n_0_126_20), .A1 (n_0_126_7), .A2 (n_0_126_9), .A3 (n_0_126_11));
NAND2_X1 i_0_126_20 (.ZN (n_0_126_19), .A1 (n_0_126_30), .A2 (\mem[5][8] ));
INV_X1 i_0_126_19 (.ZN (n_0_126_18), .A (sps__n112));
NAND4_X1 i_0_126_18 (.ZN (n_0_126_17), .A1 (n_0_126_18), .A2 (sps__n3), .A3 (sps__n122), .A4 (sps__n99));
INV_X1 i_0_126_17 (.ZN (n_0_126_16), .A (sps__n19));
INV_X1 i_0_126_16 (.ZN (n_0_126_15), .A (sps__n81));
INV_X1 i_0_126_15 (.ZN (n_0_126_14), .A (sps__n105));
NAND3_X1 i_0_126_14 (.ZN (n_0_126_13), .A1 (n_0_126_16), .A2 (n_0_126_15), .A3 (n_0_126_14));
INV_X1 i_0_126_13 (.ZN (n_0_126_12), .A (sps__n62));
INV_X1 i_0_126_12 (.ZN (n_0_126_11), .A (sps__n75));
INV_X1 i_0_126_11 (.ZN (n_0_126_10), .A (sps__n9));
INV_X1 i_0_126_10 (.ZN (n_0_126_9), .A (sps__n15));
INV_X1 i_0_126_9 (.ZN (n_0_126_8), .A (sps__n86));
INV_X1 i_0_126_8 (.ZN (n_0_126_7), .A (sps__n34));
INV_X1 i_0_126_7 (.ZN (n_0_126_6), .A (sps__n92));
INV_X1 i_0_126_6 (.ZN (n_0_126_5), .A (sps__n67));
INV_X1 i_0_126_5 (.ZN (n_0_126_4), .A (sps__n28));
INV_X1 i_0_126_4 (.ZN (n_0_126_3), .A (sps__n43));
INV_X1 i_0_126_3 (.ZN (n_0_126_2), .A (sps__n50));
INV_X1 i_0_126_2 (.ZN (n_0_126_1), .A (sps__n55));
NAND4_X1 i_0_126_1 (.ZN (n_0_126_0), .A1 (n_0_126_26), .A2 (n_0_126_25), .A3 (n_0_126_24), .A4 (data[8]));
NAND2_X1 i_0_126_0 (.ZN (n_0_115), .A1 (n_0_126_19), .A2 (n_0_126_0));
NAND3_X1 i_0_109_31 (.ZN (n_0_109_30), .A1 (n_0_109_27), .A2 (n_0_109_28), .A3 (n_0_109_29));
NOR2_X1 i_0_109_30 (.ZN (n_0_109_29), .A1 (n_0_109_13), .A2 (n_0_109_23));
NOR2_X1 i_0_109_29 (.ZN (n_0_109_28), .A1 (n_0_109_22), .A2 (n_0_109_21));
NOR2_X1 i_0_109_28 (.ZN (n_0_109_27), .A1 (n_0_109_17), .A2 (n_0_109_20));
NOR2_X1 i_0_109_27 (.ZN (n_0_109_26), .A1 (n_0_109_17), .A2 (n_0_109_13));
NOR2_X1 i_0_109_26 (.ZN (n_0_109_25), .A1 (n_0_109_20), .A2 (n_0_109_21));
NOR2_X1 i_0_109_25 (.ZN (n_0_109_24), .A1 (n_0_109_22), .A2 (n_0_109_23));
NAND3_X1 i_0_109_24 (.ZN (n_0_109_23), .A1 (n_0_109_4), .A2 (n_0_109_2), .A3 (n_0_109_6));
NAND3_X1 i_0_109_23 (.ZN (n_0_109_22), .A1 (n_0_109_1), .A2 (n_0_109_3), .A3 (n_0_109_5));
NAND3_X1 i_0_109_22 (.ZN (n_0_109_21), .A1 (n_0_109_10), .A2 (n_0_109_8), .A3 (n_0_109_12));
NAND3_X1 i_0_109_21 (.ZN (n_0_109_20), .A1 (n_0_109_7), .A2 (n_0_109_9), .A3 (n_0_109_11));
NAND2_X1 i_0_109_20 (.ZN (n_0_109_19), .A1 (n_0_109_30), .A2 (\mem[6][8] ));
INV_X1 i_0_109_19 (.ZN (n_0_109_18), .A (sps__n99));
NAND4_X1 i_0_109_18 (.ZN (n_0_109_17), .A1 (n_0_109_18), .A2 (sps__n3), .A3 (sps__n122), .A4 (sps__n112));
INV_X1 i_0_109_17 (.ZN (n_0_109_16), .A (sps__n19));
INV_X1 i_0_109_16 (.ZN (n_0_109_15), .A (sps__n81));
INV_X1 i_0_109_15 (.ZN (n_0_109_14), .A (sps__n104));
NAND3_X1 i_0_109_14 (.ZN (n_0_109_13), .A1 (n_0_109_16), .A2 (n_0_109_15), .A3 (n_0_109_14));
INV_X1 i_0_109_13 (.ZN (n_0_109_12), .A (sps__n63));
INV_X1 i_0_109_12 (.ZN (n_0_109_11), .A (sps__n75));
INV_X1 i_0_109_11 (.ZN (n_0_109_10), .A (sps__n8));
INV_X1 i_0_109_10 (.ZN (n_0_109_9), .A (sps__n15));
INV_X1 i_0_109_9 (.ZN (n_0_109_8), .A (sps__n87));
INV_X1 i_0_109_8 (.ZN (n_0_109_7), .A (sps__n34));
INV_X1 i_0_109_7 (.ZN (n_0_109_6), .A (sps__n91));
INV_X1 i_0_109_6 (.ZN (n_0_109_5), .A (sps__n67));
INV_X1 i_0_109_5 (.ZN (n_0_109_4), .A (sps__n26));
INV_X1 i_0_109_4 (.ZN (n_0_109_3), .A (sps__n43));
INV_X1 i_0_109_3 (.ZN (n_0_109_2), .A (sps__n50));
INV_X1 i_0_109_2 (.ZN (n_0_109_1), .A (sps__n57));
NAND4_X1 i_0_109_1 (.ZN (n_0_109_0), .A1 (n_0_109_26), .A2 (n_0_109_25), .A3 (n_0_109_24), .A4 (data[8]));
NAND2_X1 i_0_109_0 (.ZN (n_0_114), .A1 (n_0_109_19), .A2 (n_0_109_0));
NAND3_X1 i_0_92_27 (.ZN (n_0_92_26), .A1 (n_0_92_23), .A2 (n_0_92_24), .A3 (n_0_92_25));
NOR2_X1 i_0_92_26 (.ZN (n_0_92_25), .A1 (n_0_92_17), .A2 (n_0_92_13));
NOR2_X1 i_0_92_25 (.ZN (n_0_92_24), .A1 (n_0_92_19), .A2 (n_0_92_20));
NOR2_X1 i_0_92_24 (.ZN (n_0_92_23), .A1 (n_0_92_21), .A2 (n_0_92_22));
NAND3_X1 i_0_92_23 (.ZN (n_0_92_22), .A1 (n_0_92_4), .A2 (n_0_92_2), .A3 (n_0_92_6));
NAND3_X1 i_0_92_22 (.ZN (n_0_92_21), .A1 (n_0_92_1), .A2 (n_0_92_3), .A3 (n_0_92_5));
NAND3_X1 i_0_92_21 (.ZN (n_0_92_20), .A1 (n_0_92_10), .A2 (n_0_92_8), .A3 (n_0_92_12));
NAND3_X1 i_0_92_20 (.ZN (n_0_92_19), .A1 (n_0_92_7), .A2 (n_0_92_9), .A3 (n_0_92_11));
NAND2_X1 i_0_92_19 (.ZN (n_0_92_18), .A1 (n_0_92_26), .A2 (\mem[7][8] ));
NAND4_X1 i_0_92_18 (.ZN (n_0_92_17), .A1 (sps__n3), .A2 (sps__n122), .A3 (sps__n112), .A4 (sps__n99));
INV_X1 i_0_92_17 (.ZN (n_0_92_16), .A (sps__n19));
INV_X1 i_0_92_16 (.ZN (n_0_92_15), .A (sps__n81));
INV_X1 i_0_92_15 (.ZN (n_0_92_14), .A (sps__n105));
NAND3_X1 i_0_92_14 (.ZN (n_0_92_13), .A1 (n_0_92_16), .A2 (n_0_92_15), .A3 (n_0_92_14));
INV_X1 i_0_92_13 (.ZN (n_0_92_12), .A (sps__n62));
INV_X1 i_0_92_12 (.ZN (n_0_92_11), .A (sps__n75));
INV_X1 i_0_92_11 (.ZN (n_0_92_10), .A (sps__n9));
INV_X1 i_0_92_10 (.ZN (n_0_92_9), .A (sps__n15));
INV_X1 i_0_92_9 (.ZN (n_0_92_8), .A (sps__n86));
INV_X1 i_0_92_8 (.ZN (n_0_92_7), .A (sps__n34));
INV_X1 i_0_92_7 (.ZN (n_0_92_6), .A (sps__n92));
INV_X1 i_0_92_6 (.ZN (n_0_92_5), .A (address[6]));
INV_X1 i_0_92_5 (.ZN (n_0_92_4), .A (sps__n28));
INV_X1 i_0_92_4 (.ZN (n_0_92_3), .A (sps__n43));
INV_X1 i_0_92_3 (.ZN (n_0_92_2), .A (sps__n50));
INV_X1 i_0_92_2 (.ZN (n_0_92_1), .A (sps__n55));
NAND4_X1 i_0_92_1 (.ZN (n_0_92_0), .A1 (n_0_92_25), .A2 (n_0_92_24), .A3 (n_0_92_23), .A4 (data[8]));
NAND2_X1 i_0_92_0 (.ZN (n_0_113), .A1 (n_0_92_18), .A2 (n_0_92_0));
NAND3_X1 i_0_75_35 (.ZN (n_0_112), .A1 (n_0_75_32), .A2 (n_0_75_33), .A3 (n_0_75_34));
NAND2_X1 i_0_75_34 (.ZN (n_0_75_34), .A1 (n_0_75_23), .A2 (\mem[8][8] ));
NAND3_X1 i_0_75_29 (.ZN (n_0_75_33), .A1 (n_0_75_26), .A2 (n_0_75_31), .A3 (n_0_75_28));
NAND2_X1 i_0_75_28 (.ZN (n_0_75_32), .A1 (n_0_75_27), .A2 (\mem[8][8] ));
NOR2_X1 i_0_75_24 (.ZN (n_0_75_31), .A1 (n_0_75_18), .A2 (n_0_75_0));
INV_X1 i_0_75_23 (.ZN (n_0_75_30), .A (n_0_75_0));
INV_X1 i_0_75_22 (.ZN (n_0_75_29), .A (n_0_75_18));
INV_X1 i_0_75_21 (.ZN (n_0_75_28), .A (n_0_75_5));
NAND3_X1 i_0_75_20 (.ZN (n_0_75_27), .A1 (n_0_75_28), .A2 (n_0_75_30), .A3 (n_0_75_9));
NOR2_X1 i_0_75_19 (.ZN (n_0_75_26), .A1 (n_0_75_14), .A2 (n_0_75_24));
INV_X1 i_0_75_18 (.ZN (n_0_75_25), .A (n_0_75_14));
NAND2_X1 i_0_75_17 (.ZN (n_0_75_24), .A1 (n_0_75_9), .A2 (data[8]));
NAND2_X1 i_0_75_16 (.ZN (n_0_75_23), .A1 (n_0_75_29), .A2 (n_0_75_25));
INV_X1 i_0_75_33 (.ZN (n_0_75_22), .A (sps__n34));
INV_X1 i_0_75_32 (.ZN (n_0_75_21), .A (sps__n9));
INV_X1 i_0_75_31 (.ZN (n_0_75_20), .A (sps__n15));
INV_X1 i_0_75_30 (.ZN (n_0_75_19), .A (sps__n51));
NAND4_X1 i_0_75_3 (.ZN (n_0_75_18), .A1 (n_0_75_22), .A2 (n_0_75_21), .A3 (n_0_75_20), .A4 (n_0_75_19));
INV_X1 i_0_75_27 (.ZN (n_0_75_17), .A (sps__n63));
INV_X1 i_0_75_26 (.ZN (n_0_75_16), .A (sps__n75));
INV_X1 i_0_75_25 (.ZN (n_0_75_15), .A (sps__n87));
NAND4_X1 i_0_75_8 (.ZN (n_0_75_14), .A1 (n_0_75_17), .A2 (n_0_75_16), .A3 (n_0_75_15), .A4 (sps__n3));
INV_X1 i_0_75_15 (.ZN (n_0_75_13), .A (sps__n122));
INV_X1 i_0_75_14 (.ZN (n_0_75_12), .A (address[1]));
INV_X1 i_0_75_13 (.ZN (n_0_75_11), .A (sps__n99));
NAND3_X1 i_0_75_12 (.ZN (n_0_75_10), .A1 (n_0_75_13), .A2 (n_0_75_12), .A3 (n_0_75_11));
INV_X1 i_0_75_11 (.ZN (n_0_75_9), .A (n_0_75_10));
INV_X1 i_0_75_10 (.ZN (n_0_75_8), .A (sps__n67));
INV_X1 i_0_75_9 (.ZN (n_0_75_7), .A (sps__n19));
INV_X1 i_0_75_7 (.ZN (n_0_75_6), .A (sps__n81));
NAND4_X1 i_0_75_6 (.ZN (n_0_75_5), .A1 (n_0_75_8), .A2 (n_0_75_7), .A3 (n_0_75_6), .A4 (sps__n105));
INV_X1 i_0_75_5 (.ZN (n_0_75_4), .A (sps__n55));
INV_X1 i_0_75_4 (.ZN (n_0_75_3), .A (sps__n28));
INV_X1 i_0_75_2 (.ZN (n_0_75_2), .A (sps__n43));
INV_X1 i_0_75_1 (.ZN (n_0_75_1), .A (sps__n92));
NAND4_X1 i_0_75_0 (.ZN (n_0_75_0), .A1 (n_0_75_4), .A2 (n_0_75_3), .A3 (n_0_75_2), .A4 (n_0_75_1));
NOR2_X1 i_0_58_34 (.ZN (n_0_58_33), .A1 (n_0_58_19), .A2 (n_0_58_0));
INV_X1 i_0_58_33 (.ZN (n_0_58_32), .A (n_0_58_0));
INV_X1 i_0_58_28 (.ZN (n_0_58_31), .A (n_0_58_19));
NAND2_X1 i_0_58_27 (.ZN (n_0_58_30), .A1 (n_0_58_29), .A2 (\mem[9][8] ));
NAND3_X1 i_0_58_23 (.ZN (n_0_58_29), .A1 (n_0_58_5), .A2 (n_0_58_32), .A3 (n_0_58_10));
NAND3_X1 i_0_58_22 (.ZN (n_0_58_28), .A1 (n_0_58_27), .A2 (n_0_58_33), .A3 (n_0_58_14));
NOR2_X1 i_0_58_21 (.ZN (n_0_58_27), .A1 (n_0_58_6), .A2 (n_0_58_26));
NAND2_X1 i_0_58_20 (.ZN (n_0_58_26), .A1 (n_0_58_10), .A2 (data[8]));
NAND2_X1 i_0_58_19 (.ZN (n_0_58_25), .A1 (n_0_58_31), .A2 (n_0_58_14));
NAND3_X1 i_0_58_18 (.ZN (n_0_111), .A1 (n_0_58_28), .A2 (n_0_58_30), .A3 (n_0_58_24));
NAND2_X1 i_0_58_17 (.ZN (n_0_58_24), .A1 (n_0_58_25), .A2 (\mem[9][8] ));
INV_X1 i_0_58_32 (.ZN (n_0_58_23), .A (sps__n34));
INV_X1 i_0_58_31 (.ZN (n_0_58_22), .A (sps__n9));
INV_X1 i_0_58_30 (.ZN (n_0_58_21), .A (sps__n15));
INV_X1 i_0_58_29 (.ZN (n_0_58_20), .A (sps__n51));
NAND4_X1 i_0_58_3 (.ZN (n_0_58_19), .A1 (n_0_58_23), .A2 (n_0_58_22), .A3 (n_0_58_21), .A4 (n_0_58_20));
INV_X1 i_0_58_26 (.ZN (n_0_58_18), .A (sps__n63));
INV_X1 i_0_58_25 (.ZN (n_0_58_17), .A (sps__n75));
INV_X1 i_0_58_24 (.ZN (n_0_58_16), .A (sps__n87));
NAND4_X1 i_0_58_6 (.ZN (n_0_58_15), .A1 (n_0_58_18), .A2 (n_0_58_17), .A3 (n_0_58_16), .A4 (sps__n3));
INV_X1 i_0_58_16 (.ZN (n_0_58_14), .A (n_0_58_15));
INV_X1 i_0_58_15 (.ZN (n_0_58_13), .A (sps__n122));
INV_X1 i_0_58_14 (.ZN (n_0_58_12), .A (sps__n112));
NAND3_X1 i_0_58_13 (.ZN (n_0_58_11), .A1 (n_0_58_13), .A2 (n_0_58_12), .A3 (sps__n99));
INV_X1 i_0_58_12 (.ZN (n_0_58_10), .A (n_0_58_11));
INV_X1 i_0_58_11 (.ZN (n_0_58_9), .A (sps__n67));
INV_X1 i_0_58_10 (.ZN (n_0_58_8), .A (sps__n19));
INV_X1 i_0_58_9 (.ZN (n_0_58_7), .A (sps__n81));
NAND4_X1 i_0_58_8 (.ZN (n_0_58_6), .A1 (n_0_58_9), .A2 (n_0_58_8), .A3 (n_0_58_7), .A4 (sps__n104));
INV_X1 i_0_58_7 (.ZN (n_0_58_5), .A (n_0_58_6));
INV_X1 i_0_58_5 (.ZN (n_0_58_4), .A (sps__n57));
INV_X1 i_0_58_4 (.ZN (n_0_58_3), .A (sps__n26));
INV_X1 i_0_58_2 (.ZN (n_0_58_2), .A (sps__n43));
INV_X1 i_0_58_1 (.ZN (n_0_58_1), .A (sps__n91));
NAND4_X1 i_0_58_0 (.ZN (n_0_58_0), .A1 (n_0_58_4), .A2 (n_0_58_3), .A3 (n_0_58_2), .A4 (n_0_58_1));
NOR2_X1 i_0_41_34 (.ZN (n_0_41_33), .A1 (n_0_41_19), .A2 (n_0_41_0));
INV_X1 i_0_41_33 (.ZN (n_0_41_32), .A (n_0_41_0));
INV_X1 i_0_41_28 (.ZN (n_0_41_31), .A (n_0_41_19));
NAND2_X1 i_0_41_27 (.ZN (n_0_41_30), .A1 (n_0_41_29), .A2 (\mem[10][8] ));
NAND3_X1 i_0_41_23 (.ZN (n_0_41_29), .A1 (n_0_41_5), .A2 (n_0_41_32), .A3 (n_0_41_10));
NAND3_X1 i_0_41_22 (.ZN (n_0_41_28), .A1 (n_0_41_27), .A2 (n_0_41_33), .A3 (n_0_41_14));
NOR2_X1 i_0_41_21 (.ZN (n_0_41_27), .A1 (n_0_41_6), .A2 (n_0_41_26));
NAND2_X1 i_0_41_20 (.ZN (n_0_41_26), .A1 (n_0_41_10), .A2 (data[8]));
NAND2_X1 i_0_41_19 (.ZN (n_0_41_25), .A1 (n_0_41_31), .A2 (n_0_41_14));
NAND3_X1 i_0_41_18 (.ZN (n_0_110), .A1 (n_0_41_28), .A2 (n_0_41_30), .A3 (n_0_41_24));
NAND2_X1 i_0_41_17 (.ZN (n_0_41_24), .A1 (n_0_41_25), .A2 (\mem[10][8] ));
INV_X1 i_0_41_32 (.ZN (n_0_41_23), .A (sps__n34));
INV_X1 i_0_41_31 (.ZN (n_0_41_22), .A (sps__n9));
INV_X1 i_0_41_30 (.ZN (n_0_41_21), .A (sps__n15));
INV_X1 i_0_41_29 (.ZN (n_0_41_20), .A (sps__n51));
NAND4_X1 i_0_41_3 (.ZN (n_0_41_19), .A1 (n_0_41_23), .A2 (n_0_41_22), .A3 (n_0_41_21), .A4 (n_0_41_20));
INV_X1 i_0_41_26 (.ZN (n_0_41_18), .A (sps__n63));
INV_X1 i_0_41_25 (.ZN (n_0_41_17), .A (sps__n75));
INV_X1 i_0_41_24 (.ZN (n_0_41_16), .A (sps__n87));
NAND4_X1 i_0_41_6 (.ZN (n_0_41_15), .A1 (n_0_41_18), .A2 (n_0_41_17), .A3 (n_0_41_16), .A4 (sps__n3));
INV_X1 i_0_41_16 (.ZN (n_0_41_14), .A (n_0_41_15));
INV_X1 i_0_41_15 (.ZN (n_0_41_13), .A (sps__n122));
INV_X1 i_0_41_14 (.ZN (n_0_41_12), .A (sps__n99));
NAND3_X1 i_0_41_13 (.ZN (n_0_41_11), .A1 (n_0_41_13), .A2 (n_0_41_12), .A3 (address[1]));
INV_X1 i_0_41_12 (.ZN (n_0_41_10), .A (n_0_41_11));
INV_X1 i_0_41_11 (.ZN (n_0_41_9), .A (address[6]));
INV_X1 i_0_41_10 (.ZN (n_0_41_8), .A (sps__n19));
INV_X1 i_0_41_9 (.ZN (n_0_41_7), .A (sps__n81));
NAND4_X1 i_0_41_8 (.ZN (n_0_41_6), .A1 (n_0_41_9), .A2 (n_0_41_8), .A3 (n_0_41_7), .A4 (sps__n105));
INV_X1 i_0_41_7 (.ZN (n_0_41_5), .A (n_0_41_6));
INV_X1 i_0_41_5 (.ZN (n_0_41_4), .A (sps__n55));
INV_X1 i_0_41_4 (.ZN (n_0_41_3), .A (sps__n28));
INV_X1 i_0_41_2 (.ZN (n_0_41_2), .A (sps__n43));
INV_X1 i_0_41_1 (.ZN (n_0_41_1), .A (sps__n92));
NAND4_X1 i_0_41_0 (.ZN (n_0_41_0), .A1 (n_0_41_4), .A2 (n_0_41_3), .A3 (n_0_41_2), .A4 (n_0_41_1));
NAND3_X1 i_0_24_37 (.ZN (n_0_109), .A1 (n_0_24_34), .A2 (n_0_24_35), .A3 (n_0_24_36));
NAND2_X1 i_0_24_36 (.ZN (n_0_24_36), .A1 (n_0_24_25), .A2 (\mem[0][9] ));
NAND3_X1 i_0_24_35 (.ZN (n_0_24_35), .A1 (n_0_24_27), .A2 (n_0_24_33), .A3 (n_0_24_30));
NAND2_X1 i_0_24_34 (.ZN (n_0_24_34), .A1 (n_0_24_24), .A2 (\mem[0][9] ));
NOR2_X1 i_0_24_33 (.ZN (n_0_24_33), .A1 (n_0_24_0), .A2 (n_0_24_19));
INV_X1 i_0_24_32 (.ZN (n_0_24_32), .A (n_0_24_19));
INV_X1 i_0_24_31 (.ZN (n_0_24_31), .A (n_0_24_0));
NOR2_X1 i_0_24_30 (.ZN (n_0_24_30), .A1 (n_0_24_5), .A2 (n_0_24_15));
INV_X1 i_0_24_29 (.ZN (n_0_24_29), .A (n_0_24_15));
INV_X1 i_0_24_28 (.ZN (n_0_24_28), .A (n_0_24_5));
INV_X1 i_0_24_27 (.ZN (n_0_24_27), .A (n_0_24_26));
NAND2_X1 i_0_24_26 (.ZN (n_0_24_26), .A1 (n_0_24_10), .A2 (data[9]));
NAND2_X1 i_0_24_25 (.ZN (n_0_24_25), .A1 (n_0_24_31), .A2 (n_0_24_28));
NAND3_X1 i_0_24_24 (.ZN (n_0_24_24), .A1 (n_0_24_32), .A2 (n_0_24_29), .A3 (n_0_24_10));
INV_X1 i_0_24_23 (.ZN (n_0_24_23), .A (sps__n36));
INV_X1 i_0_24_22 (.ZN (n_0_24_22), .A (sps__n7));
INV_X1 i_0_24_21 (.ZN (n_0_24_21), .A (sps__n14));
INV_X1 i_0_24_20 (.ZN (n_0_24_20), .A (sps__n51));
NAND4_X1 i_0_24_19 (.ZN (n_0_24_19), .A1 (n_0_24_23), .A2 (n_0_24_22), .A3 (n_0_24_21), .A4 (n_0_24_20));
INV_X1 i_0_24_18 (.ZN (n_0_24_18), .A (sps__n62));
INV_X1 i_0_24_17 (.ZN (n_0_24_17), .A (sps__n74));
INV_X1 i_0_24_12 (.ZN (n_0_24_16), .A (sps__n86));
NAND4_X1 i_0_24_11 (.ZN (n_0_24_15), .A1 (n_0_24_18), .A2 (n_0_24_17), .A3 (n_0_24_16), .A4 (sps__n2));
INV_X1 i_0_24_6 (.ZN (n_0_24_14), .A (sps__n123));
INV_X1 i_0_24_5 (.ZN (n_0_24_13), .A (sps__n114));
INV_X1 i_0_24_4 (.ZN (n_0_24_12), .A (sps__n98));
NAND3_X1 i_0_24_1 (.ZN (n_0_24_11), .A1 (n_0_24_14), .A2 (n_0_24_13), .A3 (n_0_24_12));
INV_X1 i_0_24_0 (.ZN (n_0_24_10), .A (n_0_24_11));
INV_X1 i_0_24_16 (.ZN (n_0_24_9), .A (sps__n68));
INV_X1 i_0_24_15 (.ZN (n_0_24_8), .A (address[5]));
INV_X1 i_0_24_14 (.ZN (n_0_24_7), .A (address[4]));
INV_X1 i_0_24_13 (.ZN (n_0_24_6), .A (sps__n103));
NAND4_X1 i_0_24_3 (.ZN (n_0_24_5), .A1 (n_0_24_9), .A2 (n_0_24_8), .A3 (n_0_24_7), .A4 (n_0_24_6));
INV_X1 i_0_24_10 (.ZN (n_0_24_4), .A (sps__n55));
INV_X1 i_0_24_9 (.ZN (n_0_24_3), .A (address[9]));
INV_X1 i_0_24_8 (.ZN (n_0_24_2), .A (sps__n42));
INV_X1 i_0_24_7 (.ZN (n_0_24_1), .A (sps__n92));
NAND4_X1 i_0_24_2 (.ZN (n_0_24_0), .A1 (n_0_24_4), .A2 (n_0_24_3), .A3 (n_0_24_2), .A4 (n_0_24_1));
NAND3_X1 i_0_118_36 (.ZN (n_0_108), .A1 (n_0_118_33), .A2 (n_0_118_34), .A3 (n_0_118_35));
NAND2_X1 i_0_118_35 (.ZN (n_0_118_35), .A1 (n_0_118_24), .A2 (\mem[1][9] ));
NAND2_X1 i_0_118_34 (.ZN (n_0_118_34), .A1 (n_0_118_23), .A2 (\mem[1][9] ));
NAND3_X1 i_0_118_33 (.ZN (n_0_118_33), .A1 (n_0_118_26), .A2 (n_0_118_32), .A3 (n_0_118_29));
NOR2_X1 i_0_118_32 (.ZN (n_0_118_32), .A1 (n_0_118_0), .A2 (n_0_118_18));
INV_X1 i_0_118_31 (.ZN (n_0_118_31), .A (n_0_118_18));
INV_X1 i_0_118_30 (.ZN (n_0_118_30), .A (n_0_118_0));
NOR2_X1 i_0_118_29 (.ZN (n_0_118_29), .A1 (n_0_118_5), .A2 (n_0_118_14));
INV_X1 i_0_118_28 (.ZN (n_0_118_28), .A (n_0_118_14));
INV_X1 i_0_118_27 (.ZN (n_0_118_27), .A (n_0_118_5));
INV_X1 i_0_118_26 (.ZN (n_0_118_26), .A (n_0_118_25));
NAND2_X1 i_0_118_25 (.ZN (n_0_118_25), .A1 (n_0_118_10), .A2 (data[9]));
NAND2_X1 i_0_118_24 (.ZN (n_0_118_24), .A1 (n_0_118_30), .A2 (n_0_118_27));
NAND3_X1 i_0_118_23 (.ZN (n_0_118_23), .A1 (n_0_118_31), .A2 (n_0_118_28), .A3 (n_0_118_10));
INV_X1 i_0_118_22 (.ZN (n_0_118_22), .A (sps__n36));
INV_X1 i_0_118_21 (.ZN (n_0_118_21), .A (sps__n7));
INV_X1 i_0_118_20 (.ZN (n_0_118_20), .A (sps__n14));
INV_X1 i_0_118_19 (.ZN (n_0_118_19), .A (sps__n51));
NAND4_X1 i_0_118_18 (.ZN (n_0_118_18), .A1 (n_0_118_22), .A2 (n_0_118_21), .A3 (n_0_118_20), .A4 (n_0_118_19));
INV_X1 i_0_118_17 (.ZN (n_0_118_17), .A (sps__n62));
INV_X1 i_0_118_12 (.ZN (n_0_118_16), .A (sps__n74));
INV_X1 i_0_118_11 (.ZN (n_0_118_15), .A (sps__n86));
NAND4_X1 i_0_118_6 (.ZN (n_0_118_14), .A1 (n_0_118_17), .A2 (n_0_118_16), .A3 (n_0_118_15), .A4 (sps__n2));
INV_X1 i_0_118_5 (.ZN (n_0_118_13), .A (sps__n123));
INV_X1 i_0_118_4 (.ZN (n_0_118_12), .A (sps__n114));
NAND3_X1 i_0_118_1 (.ZN (n_0_118_11), .A1 (n_0_118_13), .A2 (n_0_118_12), .A3 (sps__n98));
INV_X1 i_0_118_0 (.ZN (n_0_118_10), .A (n_0_118_11));
INV_X1 i_0_118_16 (.ZN (n_0_118_9), .A (sps__n68));
INV_X1 i_0_118_15 (.ZN (n_0_118_8), .A (sps__n20));
INV_X1 i_0_118_14 (.ZN (n_0_118_7), .A (address[4]));
INV_X1 i_0_118_13 (.ZN (n_0_118_6), .A (sps__n103));
NAND4_X1 i_0_118_3 (.ZN (n_0_118_5), .A1 (n_0_118_9), .A2 (n_0_118_8), .A3 (n_0_118_7), .A4 (n_0_118_6));
INV_X1 i_0_118_10 (.ZN (n_0_118_4), .A (sps__n55));
INV_X1 i_0_118_9 (.ZN (n_0_118_3), .A (address[9]));
INV_X1 i_0_118_8 (.ZN (n_0_118_2), .A (sps__n42));
INV_X1 i_0_118_7 (.ZN (n_0_118_1), .A (sps__n92));
NAND4_X1 i_0_118_2 (.ZN (n_0_118_0), .A1 (n_0_118_4), .A2 (n_0_118_3), .A3 (n_0_118_2), .A4 (n_0_118_1));
NAND3_X1 i_0_176_36 (.ZN (n_0_107), .A1 (n_0_176_33), .A2 (n_0_176_34), .A3 (n_0_176_35));
NAND2_X1 i_0_176_35 (.ZN (n_0_176_35), .A1 (n_0_176_24), .A2 (\mem[2][9] ));
NAND2_X1 i_0_176_34 (.ZN (n_0_176_34), .A1 (n_0_176_23), .A2 (\mem[2][9] ));
NAND3_X1 i_0_176_33 (.ZN (n_0_176_33), .A1 (n_0_176_26), .A2 (n_0_176_32), .A3 (n_0_176_29));
NOR2_X1 i_0_176_32 (.ZN (n_0_176_32), .A1 (n_0_176_0), .A2 (n_0_176_18));
INV_X1 i_0_176_31 (.ZN (n_0_176_31), .A (n_0_176_18));
INV_X1 i_0_176_30 (.ZN (n_0_176_30), .A (n_0_176_0));
NOR2_X1 i_0_176_29 (.ZN (n_0_176_29), .A1 (n_0_176_5), .A2 (n_0_176_14));
INV_X1 i_0_176_28 (.ZN (n_0_176_28), .A (n_0_176_14));
INV_X1 i_0_176_27 (.ZN (n_0_176_27), .A (n_0_176_5));
INV_X1 i_0_176_26 (.ZN (n_0_176_26), .A (n_0_176_25));
NAND2_X1 i_0_176_25 (.ZN (n_0_176_25), .A1 (n_0_176_10), .A2 (data[9]));
NAND2_X1 i_0_176_24 (.ZN (n_0_176_24), .A1 (n_0_176_30), .A2 (n_0_176_27));
NAND3_X1 i_0_176_23 (.ZN (n_0_176_23), .A1 (n_0_176_31), .A2 (n_0_176_28), .A3 (n_0_176_10));
INV_X1 i_0_176_22 (.ZN (n_0_176_22), .A (sps__n36));
INV_X1 i_0_176_21 (.ZN (n_0_176_21), .A (sps__n7));
INV_X1 i_0_176_20 (.ZN (n_0_176_20), .A (sps__n14));
INV_X1 i_0_176_19 (.ZN (n_0_176_19), .A (sps__n51));
NAND4_X1 i_0_176_18 (.ZN (n_0_176_18), .A1 (n_0_176_22), .A2 (n_0_176_21), .A3 (n_0_176_20), .A4 (n_0_176_19));
INV_X1 i_0_176_17 (.ZN (n_0_176_17), .A (sps__n62));
INV_X1 i_0_176_12 (.ZN (n_0_176_16), .A (sps__n74));
INV_X1 i_0_176_11 (.ZN (n_0_176_15), .A (sps__n86));
NAND4_X1 i_0_176_6 (.ZN (n_0_176_14), .A1 (n_0_176_17), .A2 (n_0_176_16), .A3 (n_0_176_15), .A4 (sps__n2));
INV_X1 i_0_176_5 (.ZN (n_0_176_13), .A (sps__n123));
INV_X1 i_0_176_4 (.ZN (n_0_176_12), .A (sps__n98));
NAND3_X1 i_0_176_1 (.ZN (n_0_176_11), .A1 (n_0_176_13), .A2 (n_0_176_12), .A3 (sps__n114));
INV_X1 i_0_176_0 (.ZN (n_0_176_10), .A (n_0_176_11));
INV_X1 i_0_176_16 (.ZN (n_0_176_9), .A (sps__n68));
INV_X1 i_0_176_15 (.ZN (n_0_176_8), .A (address[5]));
INV_X1 i_0_176_14 (.ZN (n_0_176_7), .A (address[4]));
INV_X1 i_0_176_13 (.ZN (n_0_176_6), .A (sps__n103));
NAND4_X1 i_0_176_3 (.ZN (n_0_176_5), .A1 (n_0_176_9), .A2 (n_0_176_8), .A3 (n_0_176_7), .A4 (n_0_176_6));
INV_X1 i_0_176_10 (.ZN (n_0_176_4), .A (sps__n55));
INV_X1 i_0_176_9 (.ZN (n_0_176_3), .A (address[9]));
INV_X1 i_0_176_8 (.ZN (n_0_176_2), .A (sps__n42));
INV_X1 i_0_176_7 (.ZN (n_0_176_1), .A (sps__n92));
NAND4_X1 i_0_176_2 (.ZN (n_0_176_0), .A1 (n_0_176_4), .A2 (n_0_176_3), .A3 (n_0_176_2), .A4 (n_0_176_1));
NAND3_X1 i_0_159_31 (.ZN (n_0_159_30), .A1 (n_0_159_27), .A2 (n_0_159_28), .A3 (n_0_159_29));
NOR2_X1 i_0_159_30 (.ZN (n_0_159_29), .A1 (n_0_159_13), .A2 (n_0_159_23));
NOR2_X1 i_0_159_29 (.ZN (n_0_159_28), .A1 (n_0_159_22), .A2 (n_0_159_21));
NOR2_X1 i_0_159_28 (.ZN (n_0_159_27), .A1 (n_0_159_17), .A2 (n_0_159_20));
NOR2_X1 i_0_159_27 (.ZN (n_0_159_26), .A1 (n_0_159_17), .A2 (n_0_159_13));
NOR2_X1 i_0_159_26 (.ZN (n_0_159_25), .A1 (n_0_159_20), .A2 (n_0_159_21));
NOR2_X1 i_0_159_25 (.ZN (n_0_159_24), .A1 (n_0_159_22), .A2 (n_0_159_23));
NAND3_X1 i_0_159_24 (.ZN (n_0_159_23), .A1 (n_0_159_4), .A2 (n_0_159_2), .A3 (n_0_159_6));
NAND3_X1 i_0_159_23 (.ZN (n_0_159_22), .A1 (n_0_159_1), .A2 (n_0_159_3), .A3 (n_0_159_5));
NAND3_X1 i_0_159_22 (.ZN (n_0_159_21), .A1 (n_0_159_10), .A2 (n_0_159_8), .A3 (n_0_159_12));
NAND3_X1 i_0_159_21 (.ZN (n_0_159_20), .A1 (n_0_159_7), .A2 (n_0_159_9), .A3 (n_0_159_11));
NAND2_X1 i_0_159_20 (.ZN (n_0_159_19), .A1 (n_0_159_30), .A2 (\mem[3][9] ));
INV_X1 i_0_159_19 (.ZN (n_0_159_18), .A (sps__n123));
NAND4_X1 i_0_159_18 (.ZN (n_0_159_17), .A1 (n_0_159_18), .A2 (sps__n2), .A3 (sps__n112), .A4 (sps__n98));
INV_X1 i_0_159_17 (.ZN (n_0_159_16), .A (sps__n19));
INV_X1 i_0_159_16 (.ZN (n_0_159_15), .A (sps__n81));
INV_X1 i_0_159_15 (.ZN (n_0_159_14), .A (sps__n105));
NAND3_X1 i_0_159_14 (.ZN (n_0_159_13), .A1 (n_0_159_16), .A2 (n_0_159_15), .A3 (n_0_159_14));
INV_X1 i_0_159_13 (.ZN (n_0_159_12), .A (sps__n62));
INV_X1 i_0_159_12 (.ZN (n_0_159_11), .A (sps__n74));
INV_X1 i_0_159_11 (.ZN (n_0_159_10), .A (sps__n9));
INV_X1 i_0_159_10 (.ZN (n_0_159_9), .A (sps__n15));
INV_X1 i_0_159_9 (.ZN (n_0_159_8), .A (sps__n86));
INV_X1 i_0_159_8 (.ZN (n_0_159_7), .A (sps__n36));
INV_X1 i_0_159_7 (.ZN (n_0_159_6), .A (sps__n92));
INV_X1 i_0_159_6 (.ZN (n_0_159_5), .A (sps__n68));
INV_X1 i_0_159_5 (.ZN (n_0_159_4), .A (sps__n25));
INV_X1 i_0_159_4 (.ZN (n_0_159_3), .A (sps__n42));
INV_X1 i_0_159_3 (.ZN (n_0_159_2), .A (sps__n51));
INV_X1 i_0_159_2 (.ZN (n_0_159_1), .A (sps__n55));
NAND4_X1 i_0_159_1 (.ZN (n_0_159_0), .A1 (n_0_159_26), .A2 (n_0_159_25), .A3 (n_0_159_24), .A4 (data[9]));
NAND2_X1 i_0_159_0 (.ZN (n_0_106), .A1 (n_0_159_19), .A2 (n_0_159_0));
NAND3_X1 i_0_142_36 (.ZN (n_0_105), .A1 (n_0_142_33), .A2 (n_0_142_34), .A3 (n_0_142_35));
NAND2_X1 i_0_142_35 (.ZN (n_0_142_35), .A1 (n_0_142_24), .A2 (\mem[4][9] ));
NAND2_X1 i_0_142_34 (.ZN (n_0_142_34), .A1 (n_0_142_23), .A2 (\mem[4][9] ));
NAND3_X1 i_0_142_33 (.ZN (n_0_142_33), .A1 (n_0_142_26), .A2 (n_0_142_32), .A3 (n_0_142_29));
NOR2_X1 i_0_142_32 (.ZN (n_0_142_32), .A1 (n_0_142_0), .A2 (n_0_142_18));
INV_X1 i_0_142_31 (.ZN (n_0_142_31), .A (n_0_142_18));
INV_X1 i_0_142_30 (.ZN (n_0_142_30), .A (n_0_142_0));
NOR2_X1 i_0_142_29 (.ZN (n_0_142_29), .A1 (n_0_142_5), .A2 (n_0_142_14));
INV_X1 i_0_142_28 (.ZN (n_0_142_28), .A (n_0_142_14));
INV_X1 i_0_142_27 (.ZN (n_0_142_27), .A (n_0_142_5));
INV_X1 i_0_142_26 (.ZN (n_0_142_26), .A (n_0_142_25));
NAND2_X1 i_0_142_25 (.ZN (n_0_142_25), .A1 (n_0_142_10), .A2 (data[9]));
NAND2_X1 i_0_142_24 (.ZN (n_0_142_24), .A1 (n_0_142_30), .A2 (n_0_142_27));
NAND3_X1 i_0_142_23 (.ZN (n_0_142_23), .A1 (n_0_142_31), .A2 (n_0_142_28), .A3 (n_0_142_10));
INV_X1 i_0_142_22 (.ZN (n_0_142_22), .A (sps__n36));
INV_X1 i_0_142_21 (.ZN (n_0_142_21), .A (sps__n7));
INV_X1 i_0_142_20 (.ZN (n_0_142_20), .A (sps__n14));
INV_X1 i_0_142_19 (.ZN (n_0_142_19), .A (sps__n51));
NAND4_X1 i_0_142_18 (.ZN (n_0_142_18), .A1 (n_0_142_22), .A2 (n_0_142_21), .A3 (n_0_142_20), .A4 (n_0_142_19));
INV_X1 i_0_142_17 (.ZN (n_0_142_17), .A (sps__n62));
INV_X1 i_0_142_12 (.ZN (n_0_142_16), .A (sps__n74));
INV_X1 i_0_142_11 (.ZN (n_0_142_15), .A (sps__n86));
NAND4_X1 i_0_142_6 (.ZN (n_0_142_14), .A1 (n_0_142_17), .A2 (n_0_142_16), .A3 (n_0_142_15), .A4 (sps__n2));
INV_X1 i_0_142_5 (.ZN (n_0_142_13), .A (sps__n114));
INV_X1 i_0_142_4 (.ZN (n_0_142_12), .A (sps__n98));
NAND3_X1 i_0_142_1 (.ZN (n_0_142_11), .A1 (n_0_142_13), .A2 (n_0_142_12), .A3 (sps__n123));
INV_X1 i_0_142_0 (.ZN (n_0_142_10), .A (n_0_142_11));
INV_X1 i_0_142_16 (.ZN (n_0_142_9), .A (sps__n69));
INV_X1 i_0_142_15 (.ZN (n_0_142_8), .A (sps__n20));
INV_X1 i_0_142_14 (.ZN (n_0_142_7), .A (address[4]));
INV_X1 i_0_142_13 (.ZN (n_0_142_6), .A (sps__n103));
NAND4_X1 i_0_142_3 (.ZN (n_0_142_5), .A1 (n_0_142_9), .A2 (n_0_142_8), .A3 (n_0_142_7), .A4 (n_0_142_6));
INV_X1 i_0_142_10 (.ZN (n_0_142_4), .A (sps__n55));
INV_X1 i_0_142_9 (.ZN (n_0_142_3), .A (address[9]));
INV_X1 i_0_142_8 (.ZN (n_0_142_2), .A (sps__n42));
INV_X1 i_0_142_7 (.ZN (n_0_142_1), .A (sps__n92));
NAND4_X1 i_0_142_2 (.ZN (n_0_142_0), .A1 (n_0_142_4), .A2 (n_0_142_3), .A3 (n_0_142_2), .A4 (n_0_142_1));
NAND3_X1 i_0_125_31 (.ZN (n_0_125_30), .A1 (n_0_125_27), .A2 (n_0_125_28), .A3 (n_0_125_29));
NOR2_X1 i_0_125_30 (.ZN (n_0_125_29), .A1 (n_0_125_13), .A2 (n_0_125_23));
NOR2_X1 i_0_125_29 (.ZN (n_0_125_28), .A1 (n_0_125_22), .A2 (n_0_125_21));
NOR2_X1 i_0_125_28 (.ZN (n_0_125_27), .A1 (n_0_125_17), .A2 (n_0_125_20));
NOR2_X1 i_0_125_27 (.ZN (n_0_125_26), .A1 (n_0_125_17), .A2 (n_0_125_13));
NOR2_X1 i_0_125_26 (.ZN (n_0_125_25), .A1 (n_0_125_20), .A2 (n_0_125_21));
NOR2_X1 i_0_125_25 (.ZN (n_0_125_24), .A1 (n_0_125_22), .A2 (n_0_125_23));
NAND3_X1 i_0_125_24 (.ZN (n_0_125_23), .A1 (n_0_125_4), .A2 (n_0_125_2), .A3 (n_0_125_6));
NAND3_X1 i_0_125_23 (.ZN (n_0_125_22), .A1 (n_0_125_1), .A2 (n_0_125_3), .A3 (n_0_125_5));
NAND3_X1 i_0_125_22 (.ZN (n_0_125_21), .A1 (n_0_125_10), .A2 (n_0_125_8), .A3 (n_0_125_12));
NAND3_X1 i_0_125_21 (.ZN (n_0_125_20), .A1 (n_0_125_7), .A2 (n_0_125_9), .A3 (n_0_125_11));
NAND2_X1 i_0_125_20 (.ZN (n_0_125_19), .A1 (n_0_125_30), .A2 (\mem[5][9] ));
INV_X1 i_0_125_19 (.ZN (n_0_125_18), .A (sps__n114));
NAND4_X1 i_0_125_18 (.ZN (n_0_125_17), .A1 (n_0_125_18), .A2 (sps__n2), .A3 (sps__n123), .A4 (sps__n98));
INV_X1 i_0_125_17 (.ZN (n_0_125_16), .A (sps__n20));
INV_X1 i_0_125_16 (.ZN (n_0_125_15), .A (sps__n80));
INV_X1 i_0_125_15 (.ZN (n_0_125_14), .A (sps__n103));
NAND3_X1 i_0_125_14 (.ZN (n_0_125_13), .A1 (n_0_125_16), .A2 (n_0_125_15), .A3 (n_0_125_14));
INV_X1 i_0_125_13 (.ZN (n_0_125_12), .A (sps__n62));
INV_X1 i_0_125_12 (.ZN (n_0_125_11), .A (sps__n74));
INV_X1 i_0_125_11 (.ZN (n_0_125_10), .A (sps__n9));
INV_X1 i_0_125_10 (.ZN (n_0_125_9), .A (sps__n15));
INV_X1 i_0_125_9 (.ZN (n_0_125_8), .A (sps__n86));
INV_X1 i_0_125_8 (.ZN (n_0_125_7), .A (sps__n36));
INV_X1 i_0_125_7 (.ZN (n_0_125_6), .A (sps__n92));
INV_X1 i_0_125_6 (.ZN (n_0_125_5), .A (sps__n68));
INV_X1 i_0_125_5 (.ZN (n_0_125_4), .A (address[9]));
INV_X1 i_0_125_4 (.ZN (n_0_125_3), .A (sps__n42));
INV_X1 i_0_125_3 (.ZN (n_0_125_2), .A (sps__n51));
INV_X1 i_0_125_2 (.ZN (n_0_125_1), .A (sps__n55));
NAND4_X1 i_0_125_1 (.ZN (n_0_125_0), .A1 (n_0_125_26), .A2 (n_0_125_25), .A3 (n_0_125_24), .A4 (data[9]));
NAND2_X1 i_0_125_0 (.ZN (n_0_104), .A1 (n_0_125_19), .A2 (n_0_125_0));
NAND3_X1 i_0_108_31 (.ZN (n_0_108_30), .A1 (n_0_108_27), .A2 (n_0_108_28), .A3 (n_0_108_29));
NOR2_X1 i_0_108_30 (.ZN (n_0_108_29), .A1 (n_0_108_13), .A2 (n_0_108_23));
NOR2_X1 i_0_108_29 (.ZN (n_0_108_28), .A1 (n_0_108_22), .A2 (n_0_108_21));
NOR2_X1 i_0_108_28 (.ZN (n_0_108_27), .A1 (n_0_108_17), .A2 (n_0_108_20));
NOR2_X1 i_0_108_27 (.ZN (n_0_108_26), .A1 (n_0_108_17), .A2 (n_0_108_13));
NOR2_X1 i_0_108_26 (.ZN (n_0_108_25), .A1 (n_0_108_20), .A2 (n_0_108_21));
NOR2_X1 i_0_108_25 (.ZN (n_0_108_24), .A1 (n_0_108_22), .A2 (n_0_108_23));
NAND3_X1 i_0_108_24 (.ZN (n_0_108_23), .A1 (n_0_108_4), .A2 (n_0_108_2), .A3 (n_0_108_6));
NAND3_X1 i_0_108_23 (.ZN (n_0_108_22), .A1 (n_0_108_1), .A2 (n_0_108_3), .A3 (n_0_108_5));
NAND3_X1 i_0_108_22 (.ZN (n_0_108_21), .A1 (n_0_108_10), .A2 (n_0_108_8), .A3 (n_0_108_12));
NAND3_X1 i_0_108_21 (.ZN (n_0_108_20), .A1 (n_0_108_7), .A2 (n_0_108_9), .A3 (n_0_108_11));
NAND2_X1 i_0_108_20 (.ZN (n_0_108_19), .A1 (n_0_108_30), .A2 (\mem[6][9] ));
INV_X1 i_0_108_19 (.ZN (n_0_108_18), .A (sps__n98));
NAND4_X1 i_0_108_18 (.ZN (n_0_108_17), .A1 (n_0_108_18), .A2 (sps__n2), .A3 (sps__n123), .A4 (sps__n114));
INV_X1 i_0_108_17 (.ZN (n_0_108_16), .A (sps__n20));
INV_X1 i_0_108_16 (.ZN (n_0_108_15), .A (sps__n80));
INV_X1 i_0_108_15 (.ZN (n_0_108_14), .A (sps__n103));
NAND3_X1 i_0_108_14 (.ZN (n_0_108_13), .A1 (n_0_108_16), .A2 (n_0_108_15), .A3 (n_0_108_14));
INV_X1 i_0_108_13 (.ZN (n_0_108_12), .A (sps__n62));
INV_X1 i_0_108_12 (.ZN (n_0_108_11), .A (sps__n74));
INV_X1 i_0_108_11 (.ZN (n_0_108_10), .A (sps__n9));
INV_X1 i_0_108_10 (.ZN (n_0_108_9), .A (sps__n15));
INV_X1 i_0_108_9 (.ZN (n_0_108_8), .A (sps__n86));
INV_X1 i_0_108_8 (.ZN (n_0_108_7), .A (sps__n36));
INV_X1 i_0_108_7 (.ZN (n_0_108_6), .A (sps__n92));
INV_X1 i_0_108_6 (.ZN (n_0_108_5), .A (sps__n68));
INV_X1 i_0_108_5 (.ZN (n_0_108_4), .A (sps__n28));
INV_X1 i_0_108_4 (.ZN (n_0_108_3), .A (sps__n42));
INV_X1 i_0_108_3 (.ZN (n_0_108_2), .A (sps__n51));
INV_X1 i_0_108_2 (.ZN (n_0_108_1), .A (sps__n55));
NAND4_X1 i_0_108_1 (.ZN (n_0_108_0), .A1 (n_0_108_26), .A2 (n_0_108_25), .A3 (n_0_108_24), .A4 (data[9]));
NAND2_X1 i_0_108_0 (.ZN (n_0_103), .A1 (n_0_108_19), .A2 (n_0_108_0));
NAND3_X1 i_0_91_27 (.ZN (n_0_91_26), .A1 (n_0_91_23), .A2 (n_0_91_24), .A3 (n_0_91_25));
NOR2_X1 i_0_91_26 (.ZN (n_0_91_25), .A1 (n_0_91_17), .A2 (n_0_91_13));
NOR2_X1 i_0_91_25 (.ZN (n_0_91_24), .A1 (n_0_91_19), .A2 (n_0_91_20));
NOR2_X1 i_0_91_24 (.ZN (n_0_91_23), .A1 (n_0_91_21), .A2 (n_0_91_22));
NAND3_X1 i_0_91_23 (.ZN (n_0_91_22), .A1 (n_0_91_4), .A2 (n_0_91_2), .A3 (n_0_91_6));
NAND3_X1 i_0_91_22 (.ZN (n_0_91_21), .A1 (n_0_91_1), .A2 (n_0_91_3), .A3 (n_0_91_5));
NAND3_X1 i_0_91_21 (.ZN (n_0_91_20), .A1 (n_0_91_10), .A2 (n_0_91_8), .A3 (n_0_91_12));
NAND3_X1 i_0_91_20 (.ZN (n_0_91_19), .A1 (n_0_91_7), .A2 (n_0_91_9), .A3 (n_0_91_11));
NAND2_X1 i_0_91_19 (.ZN (n_0_91_18), .A1 (n_0_91_26), .A2 (\mem[7][9] ));
NAND4_X1 i_0_91_18 (.ZN (n_0_91_17), .A1 (sps__n2), .A2 (sps__n123), .A3 (sps__n114), .A4 (sps__n98));
INV_X1 i_0_91_17 (.ZN (n_0_91_16), .A (address[5]));
INV_X1 i_0_91_16 (.ZN (n_0_91_15), .A (address[4]));
INV_X1 i_0_91_15 (.ZN (n_0_91_14), .A (sps__n103));
NAND3_X1 i_0_91_14 (.ZN (n_0_91_13), .A1 (n_0_91_16), .A2 (n_0_91_15), .A3 (n_0_91_14));
INV_X1 i_0_91_13 (.ZN (n_0_91_12), .A (sps__n62));
INV_X1 i_0_91_12 (.ZN (n_0_91_11), .A (sps__n74));
INV_X1 i_0_91_11 (.ZN (n_0_91_10), .A (sps__n7));
INV_X1 i_0_91_10 (.ZN (n_0_91_9), .A (sps__n14));
INV_X1 i_0_91_9 (.ZN (n_0_91_8), .A (sps__n86));
INV_X1 i_0_91_8 (.ZN (n_0_91_7), .A (sps__n36));
INV_X1 i_0_91_7 (.ZN (n_0_91_6), .A (sps__n92));
INV_X1 i_0_91_6 (.ZN (n_0_91_5), .A (sps__n68));
INV_X1 i_0_91_5 (.ZN (n_0_91_4), .A (sps__n25));
INV_X1 i_0_91_4 (.ZN (n_0_91_3), .A (sps__n42));
INV_X1 i_0_91_3 (.ZN (n_0_91_2), .A (sps__n51));
INV_X1 i_0_91_2 (.ZN (n_0_91_1), .A (sps__n55));
NAND4_X1 i_0_91_1 (.ZN (n_0_91_0), .A1 (n_0_91_25), .A2 (n_0_91_24), .A3 (n_0_91_23), .A4 (data[9]));
NAND2_X1 i_0_91_0 (.ZN (n_0_102), .A1 (n_0_91_18), .A2 (n_0_91_0));
NAND3_X1 i_0_74_35 (.ZN (n_0_101), .A1 (n_0_74_32), .A2 (n_0_74_33), .A3 (n_0_74_34));
NAND2_X1 i_0_74_34 (.ZN (n_0_74_34), .A1 (n_0_74_23), .A2 (\mem[8][9] ));
NAND3_X1 i_0_74_29 (.ZN (n_0_74_33), .A1 (n_0_74_26), .A2 (n_0_74_31), .A3 (n_0_74_28));
NAND2_X1 i_0_74_28 (.ZN (n_0_74_32), .A1 (n_0_74_27), .A2 (\mem[8][9] ));
NOR2_X1 i_0_74_24 (.ZN (n_0_74_31), .A1 (n_0_74_18), .A2 (n_0_74_0));
INV_X1 i_0_74_23 (.ZN (n_0_74_30), .A (n_0_74_0));
INV_X1 i_0_74_22 (.ZN (n_0_74_29), .A (n_0_74_18));
INV_X1 i_0_74_21 (.ZN (n_0_74_28), .A (n_0_74_5));
NAND3_X1 i_0_74_20 (.ZN (n_0_74_27), .A1 (n_0_74_28), .A2 (n_0_74_30), .A3 (n_0_74_9));
NOR2_X1 i_0_74_19 (.ZN (n_0_74_26), .A1 (n_0_74_14), .A2 (n_0_74_24));
INV_X1 i_0_74_18 (.ZN (n_0_74_25), .A (n_0_74_14));
NAND2_X1 i_0_74_17 (.ZN (n_0_74_24), .A1 (n_0_74_9), .A2 (data[9]));
NAND2_X1 i_0_74_16 (.ZN (n_0_74_23), .A1 (n_0_74_29), .A2 (n_0_74_25));
INV_X1 i_0_74_33 (.ZN (n_0_74_22), .A (sps__n36));
INV_X1 i_0_74_32 (.ZN (n_0_74_21), .A (sps__n7));
INV_X1 i_0_74_31 (.ZN (n_0_74_20), .A (sps__n14));
INV_X1 i_0_74_30 (.ZN (n_0_74_19), .A (sps__n51));
NAND4_X1 i_0_74_3 (.ZN (n_0_74_18), .A1 (n_0_74_22), .A2 (n_0_74_21), .A3 (n_0_74_20), .A4 (n_0_74_19));
INV_X1 i_0_74_27 (.ZN (n_0_74_17), .A (sps__n62));
INV_X1 i_0_74_26 (.ZN (n_0_74_16), .A (sps__n74));
INV_X1 i_0_74_25 (.ZN (n_0_74_15), .A (sps__n86));
NAND4_X1 i_0_74_8 (.ZN (n_0_74_14), .A1 (n_0_74_17), .A2 (n_0_74_16), .A3 (n_0_74_15), .A4 (sps__n2));
INV_X1 i_0_74_15 (.ZN (n_0_74_13), .A (sps__n123));
INV_X1 i_0_74_14 (.ZN (n_0_74_12), .A (sps__n114));
INV_X1 i_0_74_13 (.ZN (n_0_74_11), .A (sps__n98));
NAND3_X1 i_0_74_12 (.ZN (n_0_74_10), .A1 (n_0_74_13), .A2 (n_0_74_12), .A3 (n_0_74_11));
INV_X1 i_0_74_11 (.ZN (n_0_74_9), .A (n_0_74_10));
INV_X1 i_0_74_10 (.ZN (n_0_74_8), .A (sps__n68));
INV_X1 i_0_74_9 (.ZN (n_0_74_7), .A (address[5]));
INV_X1 i_0_74_7 (.ZN (n_0_74_6), .A (address[4]));
NAND4_X1 i_0_74_6 (.ZN (n_0_74_5), .A1 (n_0_74_8), .A2 (n_0_74_7), .A3 (n_0_74_6), .A4 (sps__n103));
INV_X1 i_0_74_5 (.ZN (n_0_74_4), .A (sps__n55));
INV_X1 i_0_74_4 (.ZN (n_0_74_3), .A (address[9]));
INV_X1 i_0_74_2 (.ZN (n_0_74_2), .A (sps__n42));
INV_X1 i_0_74_1 (.ZN (n_0_74_1), .A (sps__n92));
NAND4_X1 i_0_74_0 (.ZN (n_0_74_0), .A1 (n_0_74_4), .A2 (n_0_74_3), .A3 (n_0_74_2), .A4 (n_0_74_1));
NOR2_X1 i_0_57_34 (.ZN (n_0_57_33), .A1 (n_0_57_19), .A2 (n_0_57_0));
INV_X1 i_0_57_33 (.ZN (n_0_57_32), .A (n_0_57_0));
INV_X1 i_0_57_28 (.ZN (n_0_57_31), .A (n_0_57_19));
NAND2_X1 i_0_57_27 (.ZN (n_0_57_30), .A1 (n_0_57_29), .A2 (\mem[9][9] ));
NAND3_X1 i_0_57_23 (.ZN (n_0_57_29), .A1 (n_0_57_5), .A2 (n_0_57_32), .A3 (n_0_57_10));
NAND3_X1 i_0_57_22 (.ZN (n_0_57_28), .A1 (n_0_57_27), .A2 (n_0_57_33), .A3 (n_0_57_14));
NOR2_X1 i_0_57_21 (.ZN (n_0_57_27), .A1 (n_0_57_6), .A2 (n_0_57_26));
NAND2_X1 i_0_57_20 (.ZN (n_0_57_26), .A1 (n_0_57_10), .A2 (data[9]));
NAND2_X1 i_0_57_19 (.ZN (n_0_57_25), .A1 (n_0_57_31), .A2 (n_0_57_14));
NAND3_X1 i_0_57_18 (.ZN (n_0_98), .A1 (n_0_57_28), .A2 (n_0_57_30), .A3 (n_0_57_24));
NAND2_X1 i_0_57_17 (.ZN (n_0_57_24), .A1 (n_0_57_25), .A2 (\mem[9][9] ));
INV_X1 i_0_57_32 (.ZN (n_0_57_23), .A (sps__n36));
INV_X1 i_0_57_31 (.ZN (n_0_57_22), .A (sps__n9));
INV_X1 i_0_57_30 (.ZN (n_0_57_21), .A (sps__n15));
INV_X1 i_0_57_29 (.ZN (n_0_57_20), .A (sps__n51));
NAND4_X1 i_0_57_3 (.ZN (n_0_57_19), .A1 (n_0_57_23), .A2 (n_0_57_22), .A3 (n_0_57_21), .A4 (n_0_57_20));
INV_X1 i_0_57_26 (.ZN (n_0_57_18), .A (sps__n62));
INV_X1 i_0_57_25 (.ZN (n_0_57_17), .A (sps__n74));
INV_X1 i_0_57_24 (.ZN (n_0_57_16), .A (sps__n86));
NAND4_X1 i_0_57_6 (.ZN (n_0_57_15), .A1 (n_0_57_18), .A2 (n_0_57_17), .A3 (n_0_57_16), .A4 (sps__n2));
INV_X1 i_0_57_16 (.ZN (n_0_57_14), .A (n_0_57_15));
INV_X1 i_0_57_15 (.ZN (n_0_57_13), .A (sps__n123));
INV_X1 i_0_57_14 (.ZN (n_0_57_12), .A (sps__n112));
NAND3_X1 i_0_57_13 (.ZN (n_0_57_11), .A1 (n_0_57_13), .A2 (n_0_57_12), .A3 (sps__n98));
INV_X1 i_0_57_12 (.ZN (n_0_57_10), .A (n_0_57_11));
INV_X1 i_0_57_11 (.ZN (n_0_57_9), .A (sps__n68));
INV_X1 i_0_57_10 (.ZN (n_0_57_8), .A (sps__n19));
INV_X1 i_0_57_9 (.ZN (n_0_57_7), .A (sps__n81));
NAND4_X1 i_0_57_8 (.ZN (n_0_57_6), .A1 (n_0_57_9), .A2 (n_0_57_8), .A3 (n_0_57_7), .A4 (sps__n105));
INV_X1 i_0_57_7 (.ZN (n_0_57_5), .A (n_0_57_6));
INV_X1 i_0_57_5 (.ZN (n_0_57_4), .A (sps__n55));
INV_X1 i_0_57_4 (.ZN (n_0_57_3), .A (sps__n28));
INV_X1 i_0_57_2 (.ZN (n_0_57_2), .A (sps__n43));
INV_X1 i_0_57_1 (.ZN (n_0_57_1), .A (sps__n92));
NAND4_X1 i_0_57_0 (.ZN (n_0_57_0), .A1 (n_0_57_4), .A2 (n_0_57_3), .A3 (n_0_57_2), .A4 (n_0_57_1));
NOR2_X1 i_0_40_34 (.ZN (n_0_40_33), .A1 (n_0_40_19), .A2 (n_0_40_0));
INV_X1 i_0_40_33 (.ZN (n_0_40_32), .A (n_0_40_0));
INV_X1 i_0_40_28 (.ZN (n_0_40_31), .A (n_0_40_19));
NAND2_X1 i_0_40_27 (.ZN (n_0_40_30), .A1 (n_0_40_29), .A2 (\mem[10][9] ));
NAND3_X1 i_0_40_23 (.ZN (n_0_40_29), .A1 (n_0_40_5), .A2 (n_0_40_32), .A3 (n_0_40_10));
NAND3_X1 i_0_40_22 (.ZN (n_0_40_28), .A1 (n_0_40_27), .A2 (n_0_40_33), .A3 (n_0_40_14));
NOR2_X1 i_0_40_21 (.ZN (n_0_40_27), .A1 (n_0_40_6), .A2 (n_0_40_26));
NAND2_X1 i_0_40_20 (.ZN (n_0_40_26), .A1 (n_0_40_10), .A2 (data[9]));
NAND2_X1 i_0_40_19 (.ZN (n_0_40_25), .A1 (n_0_40_31), .A2 (n_0_40_14));
NAND3_X1 i_0_40_18 (.ZN (n_0_97), .A1 (n_0_40_28), .A2 (n_0_40_30), .A3 (n_0_40_24));
NAND2_X1 i_0_40_17 (.ZN (n_0_40_24), .A1 (n_0_40_25), .A2 (\mem[10][9] ));
INV_X1 i_0_40_32 (.ZN (n_0_40_23), .A (sps__n36));
INV_X1 i_0_40_31 (.ZN (n_0_40_22), .A (sps__n9));
INV_X1 i_0_40_30 (.ZN (n_0_40_21), .A (sps__n15));
INV_X1 i_0_40_29 (.ZN (n_0_40_20), .A (sps__n51));
NAND4_X1 i_0_40_3 (.ZN (n_0_40_19), .A1 (n_0_40_23), .A2 (n_0_40_22), .A3 (n_0_40_21), .A4 (n_0_40_20));
INV_X1 i_0_40_26 (.ZN (n_0_40_18), .A (sps__n62));
INV_X1 i_0_40_25 (.ZN (n_0_40_17), .A (sps__n74));
INV_X1 i_0_40_24 (.ZN (n_0_40_16), .A (sps__n86));
NAND4_X1 i_0_40_6 (.ZN (n_0_40_15), .A1 (n_0_40_18), .A2 (n_0_40_17), .A3 (n_0_40_16), .A4 (sps__n2));
INV_X1 i_0_40_16 (.ZN (n_0_40_14), .A (n_0_40_15));
INV_X1 i_0_40_15 (.ZN (n_0_40_13), .A (sps__n123));
INV_X1 i_0_40_14 (.ZN (n_0_40_12), .A (sps__n98));
NAND3_X1 i_0_40_13 (.ZN (n_0_40_11), .A1 (n_0_40_13), .A2 (n_0_40_12), .A3 (sps__n112));
INV_X1 i_0_40_12 (.ZN (n_0_40_10), .A (n_0_40_11));
INV_X1 i_0_40_11 (.ZN (n_0_40_9), .A (sps__n68));
INV_X1 i_0_40_10 (.ZN (n_0_40_8), .A (sps__n19));
INV_X1 i_0_40_9 (.ZN (n_0_40_7), .A (sps__n81));
NAND4_X1 i_0_40_8 (.ZN (n_0_40_6), .A1 (n_0_40_9), .A2 (n_0_40_8), .A3 (n_0_40_7), .A4 (sps__n105));
INV_X1 i_0_40_7 (.ZN (n_0_40_5), .A (n_0_40_6));
INV_X1 i_0_40_5 (.ZN (n_0_40_4), .A (sps__n55));
INV_X1 i_0_40_4 (.ZN (n_0_40_3), .A (sps__n28));
INV_X1 i_0_40_2 (.ZN (n_0_40_2), .A (sps__n42));
INV_X1 i_0_40_1 (.ZN (n_0_40_1), .A (sps__n92));
NAND4_X1 i_0_40_0 (.ZN (n_0_40_0), .A1 (n_0_40_4), .A2 (n_0_40_3), .A3 (n_0_40_2), .A4 (n_0_40_1));
NAND3_X1 i_0_23_37 (.ZN (n_0_96), .A1 (n_0_23_34), .A2 (n_0_23_35), .A3 (n_0_23_36));
NAND2_X1 i_0_23_36 (.ZN (n_0_23_36), .A1 (n_0_23_25), .A2 (\mem[0][10] ));
NAND3_X1 i_0_23_35 (.ZN (n_0_23_35), .A1 (n_0_23_27), .A2 (n_0_23_33), .A3 (n_0_23_30));
NAND2_X1 i_0_23_34 (.ZN (n_0_23_34), .A1 (n_0_23_24), .A2 (\mem[0][10] ));
NOR2_X1 i_0_23_33 (.ZN (n_0_23_33), .A1 (n_0_23_0), .A2 (n_0_23_19));
INV_X1 i_0_23_32 (.ZN (n_0_23_32), .A (n_0_23_19));
INV_X1 i_0_23_31 (.ZN (n_0_23_31), .A (n_0_23_0));
NOR2_X1 i_0_23_30 (.ZN (n_0_23_30), .A1 (n_0_23_5), .A2 (n_0_23_15));
INV_X1 i_0_23_29 (.ZN (n_0_23_29), .A (n_0_23_15));
INV_X1 i_0_23_28 (.ZN (n_0_23_28), .A (n_0_23_5));
INV_X1 i_0_23_27 (.ZN (n_0_23_27), .A (n_0_23_26));
NAND2_X1 i_0_23_26 (.ZN (n_0_23_26), .A1 (n_0_23_10), .A2 (data[10]));
NAND2_X1 i_0_23_25 (.ZN (n_0_23_25), .A1 (n_0_23_31), .A2 (n_0_23_28));
NAND3_X1 i_0_23_24 (.ZN (n_0_23_24), .A1 (n_0_23_32), .A2 (n_0_23_29), .A3 (n_0_23_10));
INV_X1 i_0_23_23 (.ZN (n_0_23_23), .A (sps__n34));
INV_X1 i_0_23_22 (.ZN (n_0_23_22), .A (sps__n9));
INV_X1 i_0_23_21 (.ZN (n_0_23_21), .A (sps__n15));
INV_X1 i_0_23_20 (.ZN (n_0_23_20), .A (sps__n51));
NAND4_X1 i_0_23_19 (.ZN (n_0_23_19), .A1 (n_0_23_23), .A2 (n_0_23_22), .A3 (n_0_23_21), .A4 (n_0_23_20));
INV_X1 i_0_23_18 (.ZN (n_0_23_18), .A (sps__n62));
INV_X1 i_0_23_17 (.ZN (n_0_23_17), .A (sps__n75));
INV_X1 i_0_23_12 (.ZN (n_0_23_16), .A (sps__n86));
NAND4_X1 i_0_23_11 (.ZN (n_0_23_15), .A1 (n_0_23_18), .A2 (n_0_23_17), .A3 (n_0_23_16), .A4 (sps__n3));
INV_X1 i_0_23_6 (.ZN (n_0_23_14), .A (sps__n122));
INV_X1 i_0_23_5 (.ZN (n_0_23_13), .A (sps__n112));
INV_X1 i_0_23_4 (.ZN (n_0_23_12), .A (sps__n99));
NAND3_X1 i_0_23_1 (.ZN (n_0_23_11), .A1 (n_0_23_14), .A2 (n_0_23_13), .A3 (n_0_23_12));
INV_X1 i_0_23_0 (.ZN (n_0_23_10), .A (n_0_23_11));
INV_X1 i_0_23_16 (.ZN (n_0_23_9), .A (sps__n67));
INV_X1 i_0_23_15 (.ZN (n_0_23_8), .A (sps__n19));
INV_X1 i_0_23_14 (.ZN (n_0_23_7), .A (sps__n81));
INV_X1 i_0_23_13 (.ZN (n_0_23_6), .A (sps__n105));
NAND4_X1 i_0_23_3 (.ZN (n_0_23_5), .A1 (n_0_23_9), .A2 (n_0_23_8), .A3 (n_0_23_7), .A4 (n_0_23_6));
INV_X1 i_0_23_10 (.ZN (n_0_23_4), .A (sps__n55));
INV_X1 i_0_23_9 (.ZN (n_0_23_3), .A (sps__n25));
INV_X1 i_0_23_8 (.ZN (n_0_23_2), .A (sps__n42));
INV_X1 i_0_23_7 (.ZN (n_0_23_1), .A (sps__n92));
NAND4_X1 i_0_23_2 (.ZN (n_0_23_0), .A1 (n_0_23_4), .A2 (n_0_23_3), .A3 (n_0_23_2), .A4 (n_0_23_1));
NAND3_X1 i_0_101_36 (.ZN (n_0_95), .A1 (n_0_101_33), .A2 (n_0_101_34), .A3 (n_0_101_35));
NAND2_X1 i_0_101_35 (.ZN (n_0_101_35), .A1 (n_0_101_24), .A2 (\mem[1][10] ));
NAND2_X1 i_0_101_34 (.ZN (n_0_101_34), .A1 (n_0_101_23), .A2 (\mem[1][10] ));
NAND3_X1 i_0_101_33 (.ZN (n_0_101_33), .A1 (n_0_101_26), .A2 (n_0_101_32), .A3 (n_0_101_29));
NOR2_X1 i_0_101_32 (.ZN (n_0_101_32), .A1 (n_0_101_0), .A2 (n_0_101_18));
INV_X1 i_0_101_31 (.ZN (n_0_101_31), .A (n_0_101_18));
INV_X1 i_0_101_30 (.ZN (n_0_101_30), .A (n_0_101_0));
NOR2_X1 i_0_101_29 (.ZN (n_0_101_29), .A1 (n_0_101_5), .A2 (n_0_101_14));
INV_X1 i_0_101_28 (.ZN (n_0_101_28), .A (n_0_101_14));
INV_X1 i_0_101_27 (.ZN (n_0_101_27), .A (n_0_101_5));
INV_X1 i_0_101_26 (.ZN (n_0_101_26), .A (n_0_101_25));
NAND2_X1 i_0_101_25 (.ZN (n_0_101_25), .A1 (n_0_101_10), .A2 (data[10]));
NAND2_X1 i_0_101_24 (.ZN (n_0_101_24), .A1 (n_0_101_30), .A2 (n_0_101_27));
NAND3_X1 i_0_101_23 (.ZN (n_0_101_23), .A1 (n_0_101_31), .A2 (n_0_101_28), .A3 (n_0_101_10));
INV_X1 i_0_101_22 (.ZN (n_0_101_22), .A (sps__n34));
INV_X1 i_0_101_21 (.ZN (n_0_101_21), .A (sps__n9));
INV_X1 i_0_101_20 (.ZN (n_0_101_20), .A (sps__n15));
INV_X1 i_0_101_19 (.ZN (n_0_101_19), .A (sps__n51));
NAND4_X1 i_0_101_18 (.ZN (n_0_101_18), .A1 (n_0_101_22), .A2 (n_0_101_21), .A3 (n_0_101_20), .A4 (n_0_101_19));
INV_X1 i_0_101_17 (.ZN (n_0_101_17), .A (sps__n62));
INV_X1 i_0_101_12 (.ZN (n_0_101_16), .A (sps__n75));
INV_X1 i_0_101_11 (.ZN (n_0_101_15), .A (sps__n86));
NAND4_X1 i_0_101_6 (.ZN (n_0_101_14), .A1 (n_0_101_17), .A2 (n_0_101_16), .A3 (n_0_101_15), .A4 (sps__n3));
INV_X1 i_0_101_5 (.ZN (n_0_101_13), .A (sps__n122));
INV_X1 i_0_101_4 (.ZN (n_0_101_12), .A (sps__n112));
NAND3_X1 i_0_101_1 (.ZN (n_0_101_11), .A1 (n_0_101_13), .A2 (n_0_101_12), .A3 (sps__n99));
INV_X1 i_0_101_0 (.ZN (n_0_101_10), .A (n_0_101_11));
INV_X1 i_0_101_16 (.ZN (n_0_101_9), .A (sps__n67));
INV_X1 i_0_101_15 (.ZN (n_0_101_8), .A (sps__n19));
INV_X1 i_0_101_14 (.ZN (n_0_101_7), .A (sps__n81));
INV_X1 i_0_101_13 (.ZN (n_0_101_6), .A (sps__n105));
NAND4_X1 i_0_101_3 (.ZN (n_0_101_5), .A1 (n_0_101_9), .A2 (n_0_101_8), .A3 (n_0_101_7), .A4 (n_0_101_6));
INV_X1 i_0_101_10 (.ZN (n_0_101_4), .A (address[10]));
INV_X1 i_0_101_9 (.ZN (n_0_101_3), .A (sps__n25));
INV_X1 i_0_101_8 (.ZN (n_0_101_2), .A (sps__n42));
INV_X1 i_0_101_7 (.ZN (n_0_101_1), .A (sps__n92));
NAND4_X1 i_0_101_2 (.ZN (n_0_101_0), .A1 (n_0_101_4), .A2 (n_0_101_3), .A3 (n_0_101_2), .A4 (n_0_101_1));
NAND3_X1 i_0_175_36 (.ZN (n_0_94), .A1 (n_0_175_33), .A2 (n_0_175_34), .A3 (n_0_175_35));
NAND2_X1 i_0_175_35 (.ZN (n_0_175_35), .A1 (n_0_175_24), .A2 (\mem[2][10] ));
NAND2_X1 i_0_175_34 (.ZN (n_0_175_34), .A1 (n_0_175_23), .A2 (\mem[2][10] ));
NAND3_X1 i_0_175_33 (.ZN (n_0_175_33), .A1 (n_0_175_26), .A2 (n_0_175_32), .A3 (n_0_175_29));
NOR2_X1 i_0_175_32 (.ZN (n_0_175_32), .A1 (n_0_175_0), .A2 (n_0_175_18));
INV_X1 i_0_175_31 (.ZN (n_0_175_31), .A (n_0_175_18));
INV_X1 i_0_175_30 (.ZN (n_0_175_30), .A (n_0_175_0));
NOR2_X1 i_0_175_29 (.ZN (n_0_175_29), .A1 (n_0_175_5), .A2 (n_0_175_14));
INV_X1 i_0_175_28 (.ZN (n_0_175_28), .A (n_0_175_14));
INV_X1 i_0_175_27 (.ZN (n_0_175_27), .A (n_0_175_5));
INV_X1 i_0_175_26 (.ZN (n_0_175_26), .A (n_0_175_25));
NAND2_X1 i_0_175_25 (.ZN (n_0_175_25), .A1 (n_0_175_10), .A2 (data[10]));
NAND2_X1 i_0_175_24 (.ZN (n_0_175_24), .A1 (n_0_175_30), .A2 (n_0_175_27));
NAND3_X1 i_0_175_23 (.ZN (n_0_175_23), .A1 (n_0_175_31), .A2 (n_0_175_28), .A3 (n_0_175_10));
INV_X1 i_0_175_22 (.ZN (n_0_175_22), .A (sps__n34));
INV_X1 i_0_175_21 (.ZN (n_0_175_21), .A (sps__n9));
INV_X1 i_0_175_20 (.ZN (n_0_175_20), .A (sps__n15));
INV_X1 i_0_175_19 (.ZN (n_0_175_19), .A (sps__n51));
NAND4_X1 i_0_175_18 (.ZN (n_0_175_18), .A1 (n_0_175_22), .A2 (n_0_175_21), .A3 (n_0_175_20), .A4 (n_0_175_19));
INV_X1 i_0_175_17 (.ZN (n_0_175_17), .A (sps__n62));
INV_X1 i_0_175_12 (.ZN (n_0_175_16), .A (sps__n75));
INV_X1 i_0_175_11 (.ZN (n_0_175_15), .A (sps__n86));
NAND4_X1 i_0_175_6 (.ZN (n_0_175_14), .A1 (n_0_175_17), .A2 (n_0_175_16), .A3 (n_0_175_15), .A4 (sps__n3));
INV_X1 i_0_175_5 (.ZN (n_0_175_13), .A (sps__n122));
INV_X1 i_0_175_4 (.ZN (n_0_175_12), .A (sps__n99));
NAND3_X1 i_0_175_1 (.ZN (n_0_175_11), .A1 (n_0_175_13), .A2 (n_0_175_12), .A3 (sps__n112));
INV_X1 i_0_175_0 (.ZN (n_0_175_10), .A (n_0_175_11));
INV_X1 i_0_175_16 (.ZN (n_0_175_9), .A (sps__n68));
INV_X1 i_0_175_15 (.ZN (n_0_175_8), .A (sps__n19));
INV_X1 i_0_175_14 (.ZN (n_0_175_7), .A (sps__n81));
INV_X1 i_0_175_13 (.ZN (n_0_175_6), .A (sps__n105));
NAND4_X1 i_0_175_3 (.ZN (n_0_175_5), .A1 (n_0_175_9), .A2 (n_0_175_8), .A3 (n_0_175_7), .A4 (n_0_175_6));
INV_X1 i_0_175_10 (.ZN (n_0_175_4), .A (sps__n55));
INV_X1 i_0_175_9 (.ZN (n_0_175_3), .A (sps__n28));
INV_X1 i_0_175_8 (.ZN (n_0_175_2), .A (sps__n43));
INV_X1 i_0_175_7 (.ZN (n_0_175_1), .A (sps__n92));
NAND4_X1 i_0_175_2 (.ZN (n_0_175_0), .A1 (n_0_175_4), .A2 (n_0_175_3), .A3 (n_0_175_2), .A4 (n_0_175_1));
NAND3_X1 i_0_158_31 (.ZN (n_0_158_30), .A1 (n_0_158_27), .A2 (n_0_158_28), .A3 (n_0_158_29));
NOR2_X1 i_0_158_30 (.ZN (n_0_158_29), .A1 (n_0_158_13), .A2 (n_0_158_23));
NOR2_X1 i_0_158_29 (.ZN (n_0_158_28), .A1 (n_0_158_22), .A2 (n_0_158_21));
NOR2_X1 i_0_158_28 (.ZN (n_0_158_27), .A1 (n_0_158_17), .A2 (n_0_158_20));
NOR2_X1 i_0_158_27 (.ZN (n_0_158_26), .A1 (n_0_158_17), .A2 (n_0_158_13));
NOR2_X1 i_0_158_26 (.ZN (n_0_158_25), .A1 (n_0_158_20), .A2 (n_0_158_21));
NOR2_X1 i_0_158_25 (.ZN (n_0_158_24), .A1 (n_0_158_22), .A2 (n_0_158_23));
NAND3_X1 i_0_158_24 (.ZN (n_0_158_23), .A1 (n_0_158_4), .A2 (n_0_158_2), .A3 (n_0_158_6));
NAND3_X1 i_0_158_23 (.ZN (n_0_158_22), .A1 (n_0_158_1), .A2 (n_0_158_3), .A3 (n_0_158_5));
NAND3_X1 i_0_158_22 (.ZN (n_0_158_21), .A1 (n_0_158_10), .A2 (n_0_158_8), .A3 (n_0_158_12));
NAND3_X1 i_0_158_21 (.ZN (n_0_158_20), .A1 (n_0_158_7), .A2 (n_0_158_9), .A3 (n_0_158_11));
NAND2_X1 i_0_158_20 (.ZN (n_0_158_19), .A1 (n_0_158_30), .A2 (\mem[3][10] ));
INV_X1 i_0_158_19 (.ZN (n_0_158_18), .A (sps__n122));
NAND4_X1 i_0_158_18 (.ZN (n_0_158_17), .A1 (n_0_158_18), .A2 (sps__n2), .A3 (sps__n112), .A4 (sps__n99));
INV_X1 i_0_158_17 (.ZN (n_0_158_16), .A (sps__n19));
INV_X1 i_0_158_16 (.ZN (n_0_158_15), .A (sps__n81));
INV_X1 i_0_158_15 (.ZN (n_0_158_14), .A (sps__n105));
NAND3_X1 i_0_158_14 (.ZN (n_0_158_13), .A1 (n_0_158_16), .A2 (n_0_158_15), .A3 (n_0_158_14));
INV_X1 i_0_158_13 (.ZN (n_0_158_12), .A (sps__n62));
INV_X1 i_0_158_12 (.ZN (n_0_158_11), .A (sps__n75));
INV_X1 i_0_158_11 (.ZN (n_0_158_10), .A (sps__n9));
INV_X1 i_0_158_10 (.ZN (n_0_158_9), .A (sps__n15));
INV_X1 i_0_158_9 (.ZN (n_0_158_8), .A (sps__n86));
INV_X1 i_0_158_8 (.ZN (n_0_158_7), .A (address[14]));
INV_X1 i_0_158_7 (.ZN (n_0_158_6), .A (sps__n92));
INV_X1 i_0_158_6 (.ZN (n_0_158_5), .A (address[6]));
INV_X1 i_0_158_5 (.ZN (n_0_158_4), .A (sps__n25));
INV_X1 i_0_158_4 (.ZN (n_0_158_3), .A (sps__n42));
INV_X1 i_0_158_3 (.ZN (n_0_158_2), .A (sps__n51));
INV_X1 i_0_158_2 (.ZN (n_0_158_1), .A (address[10]));
NAND4_X1 i_0_158_1 (.ZN (n_0_158_0), .A1 (n_0_158_26), .A2 (n_0_158_25), .A3 (n_0_158_24), .A4 (data[10]));
NAND2_X1 i_0_158_0 (.ZN (n_0_93), .A1 (n_0_158_19), .A2 (n_0_158_0));
NAND3_X1 i_0_141_36 (.ZN (n_0_92), .A1 (n_0_141_33), .A2 (n_0_141_34), .A3 (n_0_141_35));
NAND2_X1 i_0_141_35 (.ZN (n_0_141_35), .A1 (n_0_141_24), .A2 (\mem[4][10] ));
NAND2_X1 i_0_141_34 (.ZN (n_0_141_34), .A1 (n_0_141_23), .A2 (\mem[4][10] ));
NAND3_X1 i_0_141_33 (.ZN (n_0_141_33), .A1 (n_0_141_26), .A2 (n_0_141_32), .A3 (n_0_141_29));
NOR2_X1 i_0_141_32 (.ZN (n_0_141_32), .A1 (n_0_141_0), .A2 (n_0_141_18));
INV_X1 i_0_141_31 (.ZN (n_0_141_31), .A (n_0_141_18));
INV_X1 i_0_141_30 (.ZN (n_0_141_30), .A (n_0_141_0));
NOR2_X1 i_0_141_29 (.ZN (n_0_141_29), .A1 (n_0_141_5), .A2 (n_0_141_14));
INV_X1 i_0_141_28 (.ZN (n_0_141_28), .A (n_0_141_14));
INV_X1 i_0_141_27 (.ZN (n_0_141_27), .A (n_0_141_5));
INV_X1 i_0_141_26 (.ZN (n_0_141_26), .A (n_0_141_25));
NAND2_X1 i_0_141_25 (.ZN (n_0_141_25), .A1 (n_0_141_10), .A2 (data[10]));
NAND2_X1 i_0_141_24 (.ZN (n_0_141_24), .A1 (n_0_141_30), .A2 (n_0_141_27));
NAND3_X1 i_0_141_23 (.ZN (n_0_141_23), .A1 (n_0_141_31), .A2 (n_0_141_28), .A3 (n_0_141_10));
INV_X1 i_0_141_22 (.ZN (n_0_141_22), .A (sps__n34));
INV_X1 i_0_141_21 (.ZN (n_0_141_21), .A (sps__n9));
INV_X1 i_0_141_20 (.ZN (n_0_141_20), .A (sps__n15));
INV_X1 i_0_141_19 (.ZN (n_0_141_19), .A (sps__n51));
NAND4_X1 i_0_141_18 (.ZN (n_0_141_18), .A1 (n_0_141_22), .A2 (n_0_141_21), .A3 (n_0_141_20), .A4 (n_0_141_19));
INV_X1 i_0_141_17 (.ZN (n_0_141_17), .A (sps__n62));
INV_X1 i_0_141_12 (.ZN (n_0_141_16), .A (sps__n75));
INV_X1 i_0_141_11 (.ZN (n_0_141_15), .A (sps__n86));
NAND4_X1 i_0_141_6 (.ZN (n_0_141_14), .A1 (n_0_141_17), .A2 (n_0_141_16), .A3 (n_0_141_15), .A4 (sps__n3));
INV_X1 i_0_141_5 (.ZN (n_0_141_13), .A (sps__n112));
INV_X1 i_0_141_4 (.ZN (n_0_141_12), .A (sps__n99));
NAND3_X1 i_0_141_1 (.ZN (n_0_141_11), .A1 (n_0_141_13), .A2 (n_0_141_12), .A3 (sps__n122));
INV_X1 i_0_141_0 (.ZN (n_0_141_10), .A (n_0_141_11));
INV_X1 i_0_141_16 (.ZN (n_0_141_9), .A (sps__n68));
INV_X1 i_0_141_15 (.ZN (n_0_141_8), .A (sps__n19));
INV_X1 i_0_141_14 (.ZN (n_0_141_7), .A (sps__n81));
INV_X1 i_0_141_13 (.ZN (n_0_141_6), .A (sps__n105));
NAND4_X1 i_0_141_3 (.ZN (n_0_141_5), .A1 (n_0_141_9), .A2 (n_0_141_8), .A3 (n_0_141_7), .A4 (n_0_141_6));
INV_X1 i_0_141_10 (.ZN (n_0_141_4), .A (sps__n55));
INV_X1 i_0_141_9 (.ZN (n_0_141_3), .A (sps__n28));
INV_X1 i_0_141_8 (.ZN (n_0_141_2), .A (sps__n43));
INV_X1 i_0_141_7 (.ZN (n_0_141_1), .A (sps__n92));
NAND4_X1 i_0_141_2 (.ZN (n_0_141_0), .A1 (n_0_141_4), .A2 (n_0_141_3), .A3 (n_0_141_2), .A4 (n_0_141_1));
NAND3_X1 i_0_124_31 (.ZN (n_0_124_30), .A1 (n_0_124_27), .A2 (n_0_124_28), .A3 (n_0_124_29));
NOR2_X1 i_0_124_30 (.ZN (n_0_124_29), .A1 (n_0_124_13), .A2 (n_0_124_23));
NOR2_X1 i_0_124_29 (.ZN (n_0_124_28), .A1 (n_0_124_22), .A2 (n_0_124_21));
NOR2_X1 i_0_124_28 (.ZN (n_0_124_27), .A1 (n_0_124_17), .A2 (n_0_124_20));
NOR2_X1 i_0_124_27 (.ZN (n_0_124_26), .A1 (n_0_124_17), .A2 (n_0_124_13));
NOR2_X1 i_0_124_26 (.ZN (n_0_124_25), .A1 (n_0_124_20), .A2 (n_0_124_21));
NOR2_X1 i_0_124_25 (.ZN (n_0_124_24), .A1 (n_0_124_22), .A2 (n_0_124_23));
NAND3_X1 i_0_124_24 (.ZN (n_0_124_23), .A1 (n_0_124_4), .A2 (n_0_124_2), .A3 (n_0_124_6));
NAND3_X1 i_0_124_23 (.ZN (n_0_124_22), .A1 (n_0_124_1), .A2 (n_0_124_3), .A3 (n_0_124_5));
NAND3_X1 i_0_124_22 (.ZN (n_0_124_21), .A1 (n_0_124_10), .A2 (n_0_124_8), .A3 (n_0_124_12));
NAND3_X1 i_0_124_21 (.ZN (n_0_124_20), .A1 (n_0_124_7), .A2 (n_0_124_9), .A3 (n_0_124_11));
NAND2_X1 i_0_124_20 (.ZN (n_0_124_19), .A1 (n_0_124_30), .A2 (\mem[5][10] ));
INV_X1 i_0_124_19 (.ZN (n_0_124_18), .A (sps__n112));
NAND4_X1 i_0_124_18 (.ZN (n_0_124_17), .A1 (n_0_124_18), .A2 (sps__n2), .A3 (sps__n122), .A4 (sps__n99));
INV_X1 i_0_124_17 (.ZN (n_0_124_16), .A (sps__n19));
INV_X1 i_0_124_16 (.ZN (n_0_124_15), .A (sps__n81));
INV_X1 i_0_124_15 (.ZN (n_0_124_14), .A (sps__n105));
NAND3_X1 i_0_124_14 (.ZN (n_0_124_13), .A1 (n_0_124_16), .A2 (n_0_124_15), .A3 (n_0_124_14));
INV_X1 i_0_124_13 (.ZN (n_0_124_12), .A (sps__n62));
INV_X1 i_0_124_12 (.ZN (n_0_124_11), .A (sps__n75));
INV_X1 i_0_124_11 (.ZN (n_0_124_10), .A (sps__n9));
INV_X1 i_0_124_10 (.ZN (n_0_124_9), .A (sps__n15));
INV_X1 i_0_124_9 (.ZN (n_0_124_8), .A (sps__n86));
INV_X1 i_0_124_8 (.ZN (n_0_124_7), .A (address[14]));
INV_X1 i_0_124_7 (.ZN (n_0_124_6), .A (sps__n92));
INV_X1 i_0_124_6 (.ZN (n_0_124_5), .A (sps__n68));
INV_X1 i_0_124_5 (.ZN (n_0_124_4), .A (sps__n28));
INV_X1 i_0_124_4 (.ZN (n_0_124_3), .A (sps__n42));
INV_X1 i_0_124_3 (.ZN (n_0_124_2), .A (sps__n51));
INV_X1 i_0_124_2 (.ZN (n_0_124_1), .A (sps__n55));
NAND4_X1 i_0_124_1 (.ZN (n_0_124_0), .A1 (n_0_124_26), .A2 (n_0_124_25), .A3 (n_0_124_24), .A4 (data[10]));
NAND2_X1 i_0_124_0 (.ZN (n_0_91), .A1 (n_0_124_19), .A2 (n_0_124_0));
NAND3_X1 i_0_107_31 (.ZN (n_0_107_30), .A1 (n_0_107_27), .A2 (n_0_107_28), .A3 (n_0_107_29));
NOR2_X1 i_0_107_30 (.ZN (n_0_107_29), .A1 (n_0_107_13), .A2 (n_0_107_23));
NOR2_X1 i_0_107_29 (.ZN (n_0_107_28), .A1 (n_0_107_22), .A2 (n_0_107_21));
NOR2_X1 i_0_107_28 (.ZN (n_0_107_27), .A1 (n_0_107_17), .A2 (n_0_107_20));
NOR2_X1 i_0_107_27 (.ZN (n_0_107_26), .A1 (n_0_107_17), .A2 (n_0_107_13));
NOR2_X1 i_0_107_26 (.ZN (n_0_107_25), .A1 (n_0_107_20), .A2 (n_0_107_21));
NOR2_X1 i_0_107_25 (.ZN (n_0_107_24), .A1 (n_0_107_22), .A2 (n_0_107_23));
NAND3_X1 i_0_107_24 (.ZN (n_0_107_23), .A1 (n_0_107_4), .A2 (n_0_107_2), .A3 (n_0_107_6));
NAND3_X1 i_0_107_23 (.ZN (n_0_107_22), .A1 (n_0_107_1), .A2 (n_0_107_3), .A3 (n_0_107_5));
NAND3_X1 i_0_107_22 (.ZN (n_0_107_21), .A1 (n_0_107_10), .A2 (n_0_107_8), .A3 (n_0_107_12));
NAND3_X1 i_0_107_21 (.ZN (n_0_107_20), .A1 (n_0_107_7), .A2 (n_0_107_9), .A3 (n_0_107_11));
NAND2_X1 i_0_107_20 (.ZN (n_0_107_19), .A1 (n_0_107_30), .A2 (\mem[6][10] ));
INV_X1 i_0_107_19 (.ZN (n_0_107_18), .A (sps__n99));
NAND4_X1 i_0_107_18 (.ZN (n_0_107_17), .A1 (n_0_107_18), .A2 (sps__n2), .A3 (sps__n122), .A4 (sps__n112));
INV_X1 i_0_107_17 (.ZN (n_0_107_16), .A (sps__n19));
INV_X1 i_0_107_16 (.ZN (n_0_107_15), .A (sps__n81));
INV_X1 i_0_107_15 (.ZN (n_0_107_14), .A (sps__n105));
NAND3_X1 i_0_107_14 (.ZN (n_0_107_13), .A1 (n_0_107_16), .A2 (n_0_107_15), .A3 (n_0_107_14));
INV_X1 i_0_107_13 (.ZN (n_0_107_12), .A (sps__n62));
INV_X1 i_0_107_12 (.ZN (n_0_107_11), .A (sps__n75));
INV_X1 i_0_107_11 (.ZN (n_0_107_10), .A (sps__n9));
INV_X1 i_0_107_10 (.ZN (n_0_107_9), .A (sps__n15));
INV_X1 i_0_107_9 (.ZN (n_0_107_8), .A (sps__n86));
INV_X1 i_0_107_8 (.ZN (n_0_107_7), .A (address[14]));
INV_X1 i_0_107_7 (.ZN (n_0_107_6), .A (sps__n92));
INV_X1 i_0_107_6 (.ZN (n_0_107_5), .A (address[6]));
INV_X1 i_0_107_5 (.ZN (n_0_107_4), .A (sps__n25));
INV_X1 i_0_107_4 (.ZN (n_0_107_3), .A (sps__n42));
INV_X1 i_0_107_3 (.ZN (n_0_107_2), .A (sps__n51));
INV_X1 i_0_107_2 (.ZN (n_0_107_1), .A (address[10]));
NAND4_X1 i_0_107_1 (.ZN (n_0_107_0), .A1 (n_0_107_26), .A2 (n_0_107_25), .A3 (n_0_107_24), .A4 (data[10]));
NAND2_X1 i_0_107_0 (.ZN (n_0_90), .A1 (n_0_107_19), .A2 (n_0_107_0));
NAND3_X1 i_0_90_27 (.ZN (n_0_90_26), .A1 (n_0_90_23), .A2 (n_0_90_24), .A3 (n_0_90_25));
NOR2_X1 i_0_90_26 (.ZN (n_0_90_25), .A1 (n_0_90_17), .A2 (n_0_90_13));
NOR2_X1 i_0_90_25 (.ZN (n_0_90_24), .A1 (n_0_90_19), .A2 (n_0_90_20));
NOR2_X1 i_0_90_24 (.ZN (n_0_90_23), .A1 (n_0_90_21), .A2 (n_0_90_22));
NAND3_X1 i_0_90_23 (.ZN (n_0_90_22), .A1 (n_0_90_4), .A2 (n_0_90_2), .A3 (n_0_90_6));
NAND3_X1 i_0_90_22 (.ZN (n_0_90_21), .A1 (n_0_90_1), .A2 (n_0_90_3), .A3 (n_0_90_5));
NAND3_X1 i_0_90_21 (.ZN (n_0_90_20), .A1 (n_0_90_10), .A2 (n_0_90_8), .A3 (n_0_90_12));
NAND3_X1 i_0_90_20 (.ZN (n_0_90_19), .A1 (n_0_90_7), .A2 (n_0_90_9), .A3 (n_0_90_11));
NAND2_X1 i_0_90_19 (.ZN (n_0_90_18), .A1 (n_0_90_26), .A2 (\mem[7][10] ));
NAND4_X1 i_0_90_18 (.ZN (n_0_90_17), .A1 (sps__n2), .A2 (sps__n122), .A3 (sps__n112), .A4 (sps__n99));
INV_X1 i_0_90_17 (.ZN (n_0_90_16), .A (sps__n19));
INV_X1 i_0_90_16 (.ZN (n_0_90_15), .A (sps__n81));
INV_X1 i_0_90_15 (.ZN (n_0_90_14), .A (sps__n105));
NAND3_X1 i_0_90_14 (.ZN (n_0_90_13), .A1 (n_0_90_16), .A2 (n_0_90_15), .A3 (n_0_90_14));
INV_X1 i_0_90_13 (.ZN (n_0_90_12), .A (sps__n62));
INV_X1 i_0_90_12 (.ZN (n_0_90_11), .A (sps__n75));
INV_X1 i_0_90_11 (.ZN (n_0_90_10), .A (sps__n9));
INV_X1 i_0_90_10 (.ZN (n_0_90_9), .A (sps__n15));
INV_X1 i_0_90_9 (.ZN (n_0_90_8), .A (sps__n86));
INV_X1 i_0_90_8 (.ZN (n_0_90_7), .A (address[14]));
INV_X1 i_0_90_7 (.ZN (n_0_90_6), .A (sps__n92));
INV_X1 i_0_90_6 (.ZN (n_0_90_5), .A (address[6]));
INV_X1 i_0_90_5 (.ZN (n_0_90_4), .A (sps__n25));
INV_X1 i_0_90_4 (.ZN (n_0_90_3), .A (sps__n42));
INV_X1 i_0_90_3 (.ZN (n_0_90_2), .A (sps__n51));
INV_X1 i_0_90_2 (.ZN (n_0_90_1), .A (address[10]));
NAND4_X1 i_0_90_1 (.ZN (n_0_90_0), .A1 (n_0_90_25), .A2 (n_0_90_24), .A3 (n_0_90_23), .A4 (data[10]));
NAND2_X1 i_0_90_0 (.ZN (n_0_89), .A1 (n_0_90_18), .A2 (n_0_90_0));
NAND3_X1 i_0_73_35 (.ZN (n_0_88), .A1 (n_0_73_32), .A2 (n_0_73_33), .A3 (n_0_73_34));
NAND2_X1 i_0_73_34 (.ZN (n_0_73_34), .A1 (n_0_73_23), .A2 (\mem[8][10] ));
NAND3_X1 i_0_73_29 (.ZN (n_0_73_33), .A1 (n_0_73_26), .A2 (n_0_73_31), .A3 (n_0_73_28));
NAND2_X1 i_0_73_28 (.ZN (n_0_73_32), .A1 (n_0_73_27), .A2 (\mem[8][10] ));
NOR2_X1 i_0_73_24 (.ZN (n_0_73_31), .A1 (n_0_73_18), .A2 (n_0_73_0));
INV_X1 i_0_73_23 (.ZN (n_0_73_30), .A (n_0_73_0));
INV_X1 i_0_73_22 (.ZN (n_0_73_29), .A (n_0_73_18));
INV_X1 i_0_73_21 (.ZN (n_0_73_28), .A (n_0_73_5));
NAND3_X1 i_0_73_20 (.ZN (n_0_73_27), .A1 (n_0_73_28), .A2 (n_0_73_30), .A3 (n_0_73_9));
NOR2_X1 i_0_73_19 (.ZN (n_0_73_26), .A1 (n_0_73_14), .A2 (n_0_73_24));
INV_X1 i_0_73_18 (.ZN (n_0_73_25), .A (n_0_73_14));
NAND2_X1 i_0_73_17 (.ZN (n_0_73_24), .A1 (n_0_73_9), .A2 (data[10]));
NAND2_X1 i_0_73_16 (.ZN (n_0_73_23), .A1 (n_0_73_29), .A2 (n_0_73_25));
INV_X1 i_0_73_33 (.ZN (n_0_73_22), .A (address[14]));
INV_X1 i_0_73_32 (.ZN (n_0_73_21), .A (sps__n9));
INV_X1 i_0_73_31 (.ZN (n_0_73_20), .A (sps__n15));
INV_X1 i_0_73_30 (.ZN (n_0_73_19), .A (sps__n51));
NAND4_X1 i_0_73_3 (.ZN (n_0_73_18), .A1 (n_0_73_22), .A2 (n_0_73_21), .A3 (n_0_73_20), .A4 (n_0_73_19));
INV_X1 i_0_73_27 (.ZN (n_0_73_17), .A (sps__n62));
INV_X1 i_0_73_26 (.ZN (n_0_73_16), .A (sps__n75));
INV_X1 i_0_73_25 (.ZN (n_0_73_15), .A (sps__n86));
NAND4_X1 i_0_73_8 (.ZN (n_0_73_14), .A1 (n_0_73_17), .A2 (n_0_73_16), .A3 (n_0_73_15), .A4 (sps__n2));
INV_X1 i_0_73_15 (.ZN (n_0_73_13), .A (sps__n122));
INV_X1 i_0_73_14 (.ZN (n_0_73_12), .A (sps__n112));
INV_X1 i_0_73_13 (.ZN (n_0_73_11), .A (sps__n99));
NAND3_X1 i_0_73_12 (.ZN (n_0_73_10), .A1 (n_0_73_13), .A2 (n_0_73_12), .A3 (n_0_73_11));
INV_X1 i_0_73_11 (.ZN (n_0_73_9), .A (n_0_73_10));
INV_X1 i_0_73_10 (.ZN (n_0_73_8), .A (sps__n68));
INV_X1 i_0_73_9 (.ZN (n_0_73_7), .A (sps__n19));
INV_X1 i_0_73_7 (.ZN (n_0_73_6), .A (sps__n81));
NAND4_X1 i_0_73_6 (.ZN (n_0_73_5), .A1 (n_0_73_8), .A2 (n_0_73_7), .A3 (n_0_73_6), .A4 (sps__n105));
INV_X1 i_0_73_5 (.ZN (n_0_73_4), .A (sps__n55));
INV_X1 i_0_73_4 (.ZN (n_0_73_3), .A (sps__n28));
INV_X1 i_0_73_2 (.ZN (n_0_73_2), .A (sps__n43));
INV_X1 i_0_73_1 (.ZN (n_0_73_1), .A (sps__n92));
NAND4_X1 i_0_73_0 (.ZN (n_0_73_0), .A1 (n_0_73_4), .A2 (n_0_73_3), .A3 (n_0_73_2), .A4 (n_0_73_1));
NOR2_X1 i_0_56_34 (.ZN (n_0_56_33), .A1 (n_0_56_19), .A2 (n_0_56_0));
INV_X1 i_0_56_33 (.ZN (n_0_56_32), .A (n_0_56_0));
INV_X1 i_0_56_28 (.ZN (n_0_56_31), .A (n_0_56_19));
NAND2_X1 i_0_56_27 (.ZN (n_0_56_30), .A1 (n_0_56_29), .A2 (\mem[9][10] ));
NAND3_X1 i_0_56_23 (.ZN (n_0_56_29), .A1 (n_0_56_5), .A2 (n_0_56_32), .A3 (n_0_56_10));
NAND3_X1 i_0_56_22 (.ZN (n_0_56_28), .A1 (n_0_56_27), .A2 (n_0_56_33), .A3 (n_0_56_14));
NOR2_X1 i_0_56_21 (.ZN (n_0_56_27), .A1 (n_0_56_6), .A2 (n_0_56_26));
NAND2_X1 i_0_56_20 (.ZN (n_0_56_26), .A1 (n_0_56_10), .A2 (data[10]));
NAND2_X1 i_0_56_19 (.ZN (n_0_56_25), .A1 (n_0_56_31), .A2 (n_0_56_14));
NAND3_X1 i_0_56_18 (.ZN (n_0_87), .A1 (n_0_56_28), .A2 (n_0_56_30), .A3 (n_0_56_24));
NAND2_X1 i_0_56_17 (.ZN (n_0_56_24), .A1 (n_0_56_25), .A2 (\mem[9][10] ));
INV_X1 i_0_56_32 (.ZN (n_0_56_23), .A (address[14]));
INV_X1 i_0_56_31 (.ZN (n_0_56_22), .A (sps__n9));
INV_X1 i_0_56_30 (.ZN (n_0_56_21), .A (sps__n15));
INV_X1 i_0_56_29 (.ZN (n_0_56_20), .A (sps__n51));
NAND4_X1 i_0_56_3 (.ZN (n_0_56_19), .A1 (n_0_56_23), .A2 (n_0_56_22), .A3 (n_0_56_21), .A4 (n_0_56_20));
INV_X1 i_0_56_26 (.ZN (n_0_56_18), .A (sps__n62));
INV_X1 i_0_56_25 (.ZN (n_0_56_17), .A (sps__n75));
INV_X1 i_0_56_24 (.ZN (n_0_56_16), .A (sps__n86));
NAND4_X1 i_0_56_6 (.ZN (n_0_56_15), .A1 (n_0_56_18), .A2 (n_0_56_17), .A3 (n_0_56_16), .A4 (sps__n2));
INV_X1 i_0_56_16 (.ZN (n_0_56_14), .A (n_0_56_15));
INV_X1 i_0_56_15 (.ZN (n_0_56_13), .A (sps__n123));
INV_X1 i_0_56_14 (.ZN (n_0_56_12), .A (sps__n112));
NAND3_X1 i_0_56_13 (.ZN (n_0_56_11), .A1 (n_0_56_13), .A2 (n_0_56_12), .A3 (sps__n99));
INV_X1 i_0_56_12 (.ZN (n_0_56_10), .A (n_0_56_11));
INV_X1 i_0_56_11 (.ZN (n_0_56_9), .A (sps__n68));
INV_X1 i_0_56_10 (.ZN (n_0_56_8), .A (sps__n19));
INV_X1 i_0_56_9 (.ZN (n_0_56_7), .A (sps__n81));
NAND4_X1 i_0_56_8 (.ZN (n_0_56_6), .A1 (n_0_56_9), .A2 (n_0_56_8), .A3 (n_0_56_7), .A4 (sps__n105));
INV_X1 i_0_56_7 (.ZN (n_0_56_5), .A (n_0_56_6));
INV_X1 i_0_56_5 (.ZN (n_0_56_4), .A (address[10]));
INV_X1 i_0_56_4 (.ZN (n_0_56_3), .A (sps__n25));
INV_X1 i_0_56_2 (.ZN (n_0_56_2), .A (sps__n42));
INV_X1 i_0_56_1 (.ZN (n_0_56_1), .A (sps__n92));
NAND4_X1 i_0_56_0 (.ZN (n_0_56_0), .A1 (n_0_56_4), .A2 (n_0_56_3), .A3 (n_0_56_2), .A4 (n_0_56_1));
NOR2_X1 i_0_39_34 (.ZN (n_0_39_33), .A1 (n_0_39_19), .A2 (n_0_39_0));
INV_X1 i_0_39_33 (.ZN (n_0_39_32), .A (n_0_39_0));
INV_X1 i_0_39_28 (.ZN (n_0_39_31), .A (n_0_39_19));
NAND2_X1 i_0_39_27 (.ZN (n_0_39_30), .A1 (n_0_39_29), .A2 (\mem[10][10] ));
NAND3_X1 i_0_39_23 (.ZN (n_0_39_29), .A1 (n_0_39_5), .A2 (n_0_39_32), .A3 (n_0_39_10));
NAND3_X1 i_0_39_22 (.ZN (n_0_39_28), .A1 (n_0_39_27), .A2 (n_0_39_33), .A3 (n_0_39_14));
NOR2_X1 i_0_39_21 (.ZN (n_0_39_27), .A1 (n_0_39_6), .A2 (n_0_39_26));
NAND2_X1 i_0_39_20 (.ZN (n_0_39_26), .A1 (n_0_39_10), .A2 (data[10]));
NAND2_X1 i_0_39_19 (.ZN (n_0_39_25), .A1 (n_0_39_31), .A2 (n_0_39_14));
NAND3_X1 i_0_39_18 (.ZN (n_0_86), .A1 (n_0_39_28), .A2 (n_0_39_30), .A3 (n_0_39_24));
NAND2_X1 i_0_39_17 (.ZN (n_0_39_24), .A1 (n_0_39_25), .A2 (\mem[10][10] ));
INV_X1 i_0_39_32 (.ZN (n_0_39_23), .A (address[14]));
INV_X1 i_0_39_31 (.ZN (n_0_39_22), .A (sps__n9));
INV_X1 i_0_39_30 (.ZN (n_0_39_21), .A (sps__n15));
INV_X1 i_0_39_29 (.ZN (n_0_39_20), .A (sps__n51));
NAND4_X1 i_0_39_3 (.ZN (n_0_39_19), .A1 (n_0_39_23), .A2 (n_0_39_22), .A3 (n_0_39_21), .A4 (n_0_39_20));
INV_X1 i_0_39_26 (.ZN (n_0_39_18), .A (sps__n62));
INV_X1 i_0_39_25 (.ZN (n_0_39_17), .A (sps__n75));
INV_X1 i_0_39_24 (.ZN (n_0_39_16), .A (sps__n86));
NAND4_X1 i_0_39_6 (.ZN (n_0_39_15), .A1 (n_0_39_18), .A2 (n_0_39_17), .A3 (n_0_39_16), .A4 (sps__n2));
INV_X1 i_0_39_16 (.ZN (n_0_39_14), .A (n_0_39_15));
INV_X1 i_0_39_15 (.ZN (n_0_39_13), .A (sps__n123));
INV_X1 i_0_39_14 (.ZN (n_0_39_12), .A (sps__n98));
NAND3_X1 i_0_39_13 (.ZN (n_0_39_11), .A1 (n_0_39_13), .A2 (n_0_39_12), .A3 (sps__n112));
INV_X1 i_0_39_12 (.ZN (n_0_39_10), .A (n_0_39_11));
INV_X1 i_0_39_11 (.ZN (n_0_39_9), .A (sps__n68));
INV_X1 i_0_39_10 (.ZN (n_0_39_8), .A (sps__n19));
INV_X1 i_0_39_9 (.ZN (n_0_39_7), .A (sps__n81));
NAND4_X1 i_0_39_8 (.ZN (n_0_39_6), .A1 (n_0_39_9), .A2 (n_0_39_8), .A3 (n_0_39_7), .A4 (sps__n105));
INV_X1 i_0_39_7 (.ZN (n_0_39_5), .A (n_0_39_6));
INV_X1 i_0_39_5 (.ZN (n_0_39_4), .A (sps__n55));
INV_X1 i_0_39_4 (.ZN (n_0_39_3), .A (sps__n28));
INV_X1 i_0_39_2 (.ZN (n_0_39_2), .A (sps__n43));
INV_X1 i_0_39_1 (.ZN (n_0_39_1), .A (sps__n92));
NAND4_X1 i_0_39_0 (.ZN (n_0_39_0), .A1 (n_0_39_4), .A2 (n_0_39_3), .A3 (n_0_39_2), .A4 (n_0_39_1));
NAND3_X1 i_0_22_37 (.ZN (n_0_85), .A1 (n_0_22_34), .A2 (n_0_22_35), .A3 (n_0_22_36));
NAND2_X1 i_0_22_36 (.ZN (n_0_22_36), .A1 (n_0_22_25), .A2 (\mem[0][11] ));
NAND3_X1 i_0_22_35 (.ZN (n_0_22_35), .A1 (n_0_22_27), .A2 (n_0_22_33), .A3 (n_0_22_30));
NAND2_X1 i_0_22_34 (.ZN (n_0_22_34), .A1 (n_0_22_24), .A2 (\mem[0][11] ));
NOR2_X1 i_0_22_33 (.ZN (n_0_22_33), .A1 (n_0_22_0), .A2 (n_0_22_19));
INV_X1 i_0_22_32 (.ZN (n_0_22_32), .A (n_0_22_19));
INV_X1 i_0_22_31 (.ZN (n_0_22_31), .A (n_0_22_0));
NOR2_X1 i_0_22_30 (.ZN (n_0_22_30), .A1 (n_0_22_5), .A2 (n_0_22_15));
INV_X1 i_0_22_29 (.ZN (n_0_22_29), .A (n_0_22_15));
INV_X1 i_0_22_28 (.ZN (n_0_22_28), .A (n_0_22_5));
INV_X1 i_0_22_27 (.ZN (n_0_22_27), .A (n_0_22_26));
NAND2_X1 i_0_22_26 (.ZN (n_0_22_26), .A1 (n_0_22_10), .A2 (data[11]));
NAND2_X1 i_0_22_25 (.ZN (n_0_22_25), .A1 (n_0_22_31), .A2 (n_0_22_28));
NAND3_X1 i_0_22_24 (.ZN (n_0_22_24), .A1 (n_0_22_32), .A2 (n_0_22_29), .A3 (n_0_22_10));
INV_X1 i_0_22_23 (.ZN (n_0_22_23), .A (sps__n36));
INV_X1 i_0_22_22 (.ZN (n_0_22_22), .A (sps__n9));
INV_X1 i_0_22_21 (.ZN (n_0_22_21), .A (sps__n15));
INV_X1 i_0_22_20 (.ZN (n_0_22_20), .A (sps__n50));
NAND4_X1 i_0_22_19 (.ZN (n_0_22_19), .A1 (n_0_22_23), .A2 (n_0_22_22), .A3 (n_0_22_21), .A4 (n_0_22_20));
INV_X1 i_0_22_18 (.ZN (n_0_22_18), .A (sps__n62));
INV_X1 i_0_22_17 (.ZN (n_0_22_17), .A (sps__n74));
INV_X1 i_0_22_12 (.ZN (n_0_22_16), .A (sps__n86));
NAND4_X1 i_0_22_11 (.ZN (n_0_22_15), .A1 (n_0_22_18), .A2 (n_0_22_17), .A3 (n_0_22_16), .A4 (sps__n2));
INV_X1 i_0_22_6 (.ZN (n_0_22_14), .A (sps__n123));
INV_X1 i_0_22_5 (.ZN (n_0_22_13), .A (sps__n112));
INV_X1 i_0_22_4 (.ZN (n_0_22_12), .A (sps__n98));
NAND3_X1 i_0_22_1 (.ZN (n_0_22_11), .A1 (n_0_22_14), .A2 (n_0_22_13), .A3 (n_0_22_12));
INV_X1 i_0_22_0 (.ZN (n_0_22_10), .A (n_0_22_11));
INV_X1 i_0_22_16 (.ZN (n_0_22_9), .A (sps__n68));
INV_X1 i_0_22_15 (.ZN (n_0_22_8), .A (sps__n19));
INV_X1 i_0_22_14 (.ZN (n_0_22_7), .A (sps__n81));
INV_X1 i_0_22_13 (.ZN (n_0_22_6), .A (sps__n104));
NAND4_X1 i_0_22_3 (.ZN (n_0_22_5), .A1 (n_0_22_9), .A2 (n_0_22_8), .A3 (n_0_22_7), .A4 (n_0_22_6));
INV_X1 i_0_22_10 (.ZN (n_0_22_4), .A (sps__n55));
INV_X1 i_0_22_9 (.ZN (n_0_22_3), .A (sps__n28));
INV_X1 i_0_22_8 (.ZN (n_0_22_2), .A (sps__n42));
INV_X1 i_0_22_7 (.ZN (n_0_22_1), .A (sps__n92));
NAND4_X1 i_0_22_2 (.ZN (n_0_22_0), .A1 (n_0_22_4), .A2 (n_0_22_3), .A3 (n_0_22_2), .A4 (n_0_22_1));
NAND3_X1 i_0_16_36 (.ZN (n_0_84), .A1 (n_0_16_33), .A2 (n_0_16_34), .A3 (n_0_16_35));
NAND2_X1 i_0_16_35 (.ZN (n_0_16_35), .A1 (n_0_16_24), .A2 (\mem[1][11] ));
NAND2_X1 i_0_16_34 (.ZN (n_0_16_34), .A1 (n_0_16_23), .A2 (\mem[1][11] ));
NAND3_X1 i_0_16_33 (.ZN (n_0_16_33), .A1 (n_0_16_26), .A2 (n_0_16_32), .A3 (n_0_16_29));
NOR2_X1 i_0_16_32 (.ZN (n_0_16_32), .A1 (n_0_16_0), .A2 (n_0_16_18));
INV_X1 i_0_16_31 (.ZN (n_0_16_31), .A (n_0_16_18));
INV_X1 i_0_16_30 (.ZN (n_0_16_30), .A (n_0_16_0));
NOR2_X1 i_0_16_29 (.ZN (n_0_16_29), .A1 (n_0_16_5), .A2 (n_0_16_14));
INV_X1 i_0_16_28 (.ZN (n_0_16_28), .A (n_0_16_14));
INV_X1 i_0_16_27 (.ZN (n_0_16_27), .A (n_0_16_5));
INV_X1 i_0_16_26 (.ZN (n_0_16_26), .A (n_0_16_25));
NAND2_X1 i_0_16_25 (.ZN (n_0_16_25), .A1 (n_0_16_10), .A2 (data[11]));
NAND2_X1 i_0_16_24 (.ZN (n_0_16_24), .A1 (n_0_16_30), .A2 (n_0_16_27));
NAND3_X1 i_0_16_23 (.ZN (n_0_16_23), .A1 (n_0_16_31), .A2 (n_0_16_28), .A3 (n_0_16_10));
INV_X1 i_0_16_22 (.ZN (n_0_16_22), .A (sps__n35));
INV_X1 i_0_16_21 (.ZN (n_0_16_21), .A (sps__n8));
INV_X1 i_0_16_20 (.ZN (n_0_16_20), .A (sps__n13));
INV_X1 i_0_16_19 (.ZN (n_0_16_19), .A (sps__n49));
NAND4_X1 i_0_16_18 (.ZN (n_0_16_18), .A1 (n_0_16_22), .A2 (n_0_16_21), .A3 (n_0_16_20), .A4 (n_0_16_19));
INV_X1 i_0_16_17 (.ZN (n_0_16_17), .A (sps__n63));
INV_X1 i_0_16_12 (.ZN (n_0_16_16), .A (sps__n74));
INV_X1 i_0_16_11 (.ZN (n_0_16_15), .A (sps__n87));
NAND4_X1 i_0_16_6 (.ZN (n_0_16_14), .A1 (n_0_16_17), .A2 (n_0_16_16), .A3 (n_0_16_15), .A4 (sps__n1));
INV_X1 i_0_16_5 (.ZN (n_0_16_13), .A (sps__n121));
INV_X1 i_0_16_4 (.ZN (n_0_16_12), .A (sps__n112));
NAND3_X1 i_0_16_1 (.ZN (n_0_16_11), .A1 (n_0_16_13), .A2 (n_0_16_12), .A3 (sps__n97));
INV_X1 i_0_16_0 (.ZN (n_0_16_10), .A (n_0_16_11));
INV_X1 i_0_16_16 (.ZN (n_0_16_9), .A (sps__n67));
INV_X1 i_0_16_15 (.ZN (n_0_16_8), .A (sps__n21));
INV_X1 i_0_16_14 (.ZN (n_0_16_7), .A (sps__n80));
INV_X1 i_0_16_13 (.ZN (n_0_16_6), .A (sps__n106));
NAND4_X1 i_0_16_3 (.ZN (n_0_16_5), .A1 (n_0_16_9), .A2 (n_0_16_8), .A3 (n_0_16_7), .A4 (n_0_16_6));
INV_X1 i_0_16_10 (.ZN (n_0_16_4), .A (sps__n57));
INV_X1 i_0_16_9 (.ZN (n_0_16_3), .A (sps__n27));
INV_X1 i_0_16_8 (.ZN (n_0_16_2), .A (sps__n44));
INV_X1 i_0_16_7 (.ZN (n_0_16_1), .A (sps__n93));
NAND4_X1 i_0_16_2 (.ZN (n_0_16_0), .A1 (n_0_16_4), .A2 (n_0_16_3), .A3 (n_0_16_2), .A4 (n_0_16_1));
NAND3_X1 i_0_174_36 (.ZN (n_0_83), .A1 (n_0_174_33), .A2 (n_0_174_34), .A3 (n_0_174_35));
NAND2_X1 i_0_174_35 (.ZN (n_0_174_35), .A1 (n_0_174_24), .A2 (\mem[2][11] ));
NAND2_X1 i_0_174_34 (.ZN (n_0_174_34), .A1 (n_0_174_23), .A2 (\mem[2][11] ));
NAND3_X1 i_0_174_33 (.ZN (n_0_174_33), .A1 (n_0_174_26), .A2 (n_0_174_32), .A3 (n_0_174_29));
NOR2_X1 i_0_174_32 (.ZN (n_0_174_32), .A1 (n_0_174_0), .A2 (n_0_174_18));
INV_X1 i_0_174_31 (.ZN (n_0_174_31), .A (n_0_174_18));
INV_X1 i_0_174_30 (.ZN (n_0_174_30), .A (n_0_174_0));
NOR2_X1 i_0_174_29 (.ZN (n_0_174_29), .A1 (n_0_174_5), .A2 (n_0_174_14));
INV_X1 i_0_174_28 (.ZN (n_0_174_28), .A (n_0_174_14));
INV_X1 i_0_174_27 (.ZN (n_0_174_27), .A (n_0_174_5));
INV_X1 i_0_174_26 (.ZN (n_0_174_26), .A (n_0_174_25));
NAND2_X1 i_0_174_25 (.ZN (n_0_174_25), .A1 (n_0_174_10), .A2 (data[11]));
NAND2_X1 i_0_174_24 (.ZN (n_0_174_24), .A1 (n_0_174_30), .A2 (n_0_174_27));
NAND3_X1 i_0_174_23 (.ZN (n_0_174_23), .A1 (n_0_174_31), .A2 (n_0_174_28), .A3 (n_0_174_10));
INV_X1 i_0_174_22 (.ZN (n_0_174_22), .A (sps__n34));
INV_X1 i_0_174_21 (.ZN (n_0_174_21), .A (sps__n9));
INV_X1 i_0_174_20 (.ZN (n_0_174_20), .A (sps__n15));
INV_X1 i_0_174_19 (.ZN (n_0_174_19), .A (sps__n51));
NAND4_X1 i_0_174_18 (.ZN (n_0_174_18), .A1 (n_0_174_22), .A2 (n_0_174_21), .A3 (n_0_174_20), .A4 (n_0_174_19));
INV_X1 i_0_174_17 (.ZN (n_0_174_17), .A (sps__n62));
INV_X1 i_0_174_12 (.ZN (n_0_174_16), .A (sps__n74));
INV_X1 i_0_174_11 (.ZN (n_0_174_15), .A (sps__n86));
NAND4_X1 i_0_174_6 (.ZN (n_0_174_14), .A1 (n_0_174_17), .A2 (n_0_174_16), .A3 (n_0_174_15), .A4 (sps__n3));
INV_X1 i_0_174_5 (.ZN (n_0_174_13), .A (sps__n121));
INV_X1 i_0_174_4 (.ZN (n_0_174_12), .A (sps__n99));
NAND3_X1 i_0_174_1 (.ZN (n_0_174_11), .A1 (n_0_174_13), .A2 (n_0_174_12), .A3 (sps__n112));
INV_X1 i_0_174_0 (.ZN (n_0_174_10), .A (n_0_174_11));
INV_X1 i_0_174_16 (.ZN (n_0_174_9), .A (sps__n68));
INV_X1 i_0_174_15 (.ZN (n_0_174_8), .A (sps__n19));
INV_X1 i_0_174_14 (.ZN (n_0_174_7), .A (sps__n81));
INV_X1 i_0_174_13 (.ZN (n_0_174_6), .A (sps__n104));
NAND4_X1 i_0_174_3 (.ZN (n_0_174_5), .A1 (n_0_174_9), .A2 (n_0_174_8), .A3 (n_0_174_7), .A4 (n_0_174_6));
INV_X1 i_0_174_10 (.ZN (n_0_174_4), .A (sps__n55));
INV_X1 i_0_174_9 (.ZN (n_0_174_3), .A (sps__n28));
INV_X1 i_0_174_8 (.ZN (n_0_174_2), .A (sps__n43));
INV_X1 i_0_174_7 (.ZN (n_0_174_1), .A (sps__n92));
NAND4_X1 i_0_174_2 (.ZN (n_0_174_0), .A1 (n_0_174_4), .A2 (n_0_174_3), .A3 (n_0_174_2), .A4 (n_0_174_1));
NAND3_X1 i_0_157_31 (.ZN (n_0_157_30), .A1 (n_0_157_27), .A2 (n_0_157_28), .A3 (n_0_157_29));
NOR2_X1 i_0_157_30 (.ZN (n_0_157_29), .A1 (n_0_157_13), .A2 (n_0_157_23));
NOR2_X1 i_0_157_29 (.ZN (n_0_157_28), .A1 (n_0_157_22), .A2 (n_0_157_21));
NOR2_X1 i_0_157_28 (.ZN (n_0_157_27), .A1 (n_0_157_17), .A2 (n_0_157_20));
NOR2_X1 i_0_157_27 (.ZN (n_0_157_26), .A1 (n_0_157_17), .A2 (n_0_157_13));
NOR2_X1 i_0_157_26 (.ZN (n_0_157_25), .A1 (n_0_157_20), .A2 (n_0_157_21));
NOR2_X1 i_0_157_25 (.ZN (n_0_157_24), .A1 (n_0_157_22), .A2 (n_0_157_23));
NAND3_X1 i_0_157_24 (.ZN (n_0_157_23), .A1 (n_0_157_4), .A2 (n_0_157_2), .A3 (n_0_157_6));
NAND3_X1 i_0_157_23 (.ZN (n_0_157_22), .A1 (n_0_157_1), .A2 (n_0_157_3), .A3 (n_0_157_5));
NAND3_X1 i_0_157_22 (.ZN (n_0_157_21), .A1 (n_0_157_10), .A2 (n_0_157_8), .A3 (n_0_157_12));
NAND3_X1 i_0_157_21 (.ZN (n_0_157_20), .A1 (n_0_157_7), .A2 (n_0_157_9), .A3 (n_0_157_11));
NAND2_X1 i_0_157_20 (.ZN (n_0_157_19), .A1 (n_0_157_30), .A2 (\mem[3][11] ));
INV_X1 i_0_157_19 (.ZN (n_0_157_18), .A (sps__n121));
NAND4_X1 i_0_157_18 (.ZN (n_0_157_17), .A1 (n_0_157_18), .A2 (sps__n2), .A3 (sps__n114), .A4 (sps__n97));
INV_X1 i_0_157_17 (.ZN (n_0_157_16), .A (sps__n21));
INV_X1 i_0_157_16 (.ZN (n_0_157_15), .A (sps__n80));
INV_X1 i_0_157_15 (.ZN (n_0_157_14), .A (sps__n103));
NAND3_X1 i_0_157_14 (.ZN (n_0_157_13), .A1 (n_0_157_16), .A2 (n_0_157_15), .A3 (n_0_157_14));
INV_X1 i_0_157_13 (.ZN (n_0_157_12), .A (sps__n61));
INV_X1 i_0_157_12 (.ZN (n_0_157_11), .A (sps__n74));
INV_X1 i_0_157_11 (.ZN (n_0_157_10), .A (sps__n7));
INV_X1 i_0_157_10 (.ZN (n_0_157_9), .A (sps__n14));
INV_X1 i_0_157_9 (.ZN (n_0_157_8), .A (sps__n85));
INV_X1 i_0_157_8 (.ZN (n_0_157_7), .A (sps__n36));
INV_X1 i_0_157_7 (.ZN (n_0_157_6), .A (sps__n91));
INV_X1 i_0_157_6 (.ZN (n_0_157_5), .A (sps__n69));
INV_X1 i_0_157_5 (.ZN (n_0_157_4), .A (sps__n26));
INV_X1 i_0_157_4 (.ZN (n_0_157_3), .A (sps__n41));
INV_X1 i_0_157_3 (.ZN (n_0_157_2), .A (sps__n49));
INV_X1 i_0_157_2 (.ZN (n_0_157_1), .A (sps__n56));
NAND4_X1 i_0_157_1 (.ZN (n_0_157_0), .A1 (n_0_157_26), .A2 (n_0_157_25), .A3 (n_0_157_24), .A4 (data[11]));
NAND2_X1 i_0_157_0 (.ZN (n_0_82), .A1 (n_0_157_19), .A2 (n_0_157_0));
NAND3_X1 i_0_140_36 (.ZN (n_0_81), .A1 (n_0_140_33), .A2 (n_0_140_34), .A3 (n_0_140_35));
NAND2_X1 i_0_140_35 (.ZN (n_0_140_35), .A1 (n_0_140_24), .A2 (\mem[4][11] ));
NAND2_X1 i_0_140_34 (.ZN (n_0_140_34), .A1 (n_0_140_23), .A2 (\mem[4][11] ));
NAND3_X1 i_0_140_33 (.ZN (n_0_140_33), .A1 (n_0_140_26), .A2 (n_0_140_32), .A3 (n_0_140_29));
NOR2_X1 i_0_140_32 (.ZN (n_0_140_32), .A1 (n_0_140_0), .A2 (n_0_140_18));
INV_X1 i_0_140_31 (.ZN (n_0_140_31), .A (n_0_140_18));
INV_X1 i_0_140_30 (.ZN (n_0_140_30), .A (n_0_140_0));
NOR2_X1 i_0_140_29 (.ZN (n_0_140_29), .A1 (n_0_140_5), .A2 (n_0_140_14));
INV_X1 i_0_140_28 (.ZN (n_0_140_28), .A (n_0_140_14));
INV_X1 i_0_140_27 (.ZN (n_0_140_27), .A (n_0_140_5));
INV_X1 i_0_140_26 (.ZN (n_0_140_26), .A (n_0_140_25));
NAND2_X1 i_0_140_25 (.ZN (n_0_140_25), .A1 (n_0_140_10), .A2 (data[11]));
NAND2_X1 i_0_140_24 (.ZN (n_0_140_24), .A1 (n_0_140_30), .A2 (n_0_140_27));
NAND3_X1 i_0_140_23 (.ZN (n_0_140_23), .A1 (n_0_140_31), .A2 (n_0_140_28), .A3 (n_0_140_10));
INV_X1 i_0_140_22 (.ZN (n_0_140_22), .A (sps__n36));
INV_X1 i_0_140_21 (.ZN (n_0_140_21), .A (sps__n9));
INV_X1 i_0_140_20 (.ZN (n_0_140_20), .A (sps__n15));
INV_X1 i_0_140_19 (.ZN (n_0_140_19), .A (sps__n51));
NAND4_X1 i_0_140_18 (.ZN (n_0_140_18), .A1 (n_0_140_22), .A2 (n_0_140_21), .A3 (n_0_140_20), .A4 (n_0_140_19));
INV_X1 i_0_140_17 (.ZN (n_0_140_17), .A (sps__n62));
INV_X1 i_0_140_12 (.ZN (n_0_140_16), .A (sps__n74));
INV_X1 i_0_140_11 (.ZN (n_0_140_15), .A (sps__n86));
NAND4_X1 i_0_140_6 (.ZN (n_0_140_14), .A1 (n_0_140_17), .A2 (n_0_140_16), .A3 (n_0_140_15), .A4 (sps__n2));
INV_X1 i_0_140_5 (.ZN (n_0_140_13), .A (sps__n112));
INV_X1 i_0_140_4 (.ZN (n_0_140_12), .A (sps__n98));
NAND3_X1 i_0_140_1 (.ZN (n_0_140_11), .A1 (n_0_140_13), .A2 (n_0_140_12), .A3 (sps__n123));
INV_X1 i_0_140_0 (.ZN (n_0_140_10), .A (n_0_140_11));
INV_X1 i_0_140_16 (.ZN (n_0_140_9), .A (sps__n68));
INV_X1 i_0_140_15 (.ZN (n_0_140_8), .A (sps__n19));
INV_X1 i_0_140_14 (.ZN (n_0_140_7), .A (sps__n81));
INV_X1 i_0_140_13 (.ZN (n_0_140_6), .A (sps__n105));
NAND4_X1 i_0_140_3 (.ZN (n_0_140_5), .A1 (n_0_140_9), .A2 (n_0_140_8), .A3 (n_0_140_7), .A4 (n_0_140_6));
INV_X1 i_0_140_10 (.ZN (n_0_140_4), .A (sps__n55));
INV_X1 i_0_140_9 (.ZN (n_0_140_3), .A (sps__n28));
INV_X1 i_0_140_8 (.ZN (n_0_140_2), .A (sps__n43));
INV_X1 i_0_140_7 (.ZN (n_0_140_1), .A (sps__n92));
NAND4_X1 i_0_140_2 (.ZN (n_0_140_0), .A1 (n_0_140_4), .A2 (n_0_140_3), .A3 (n_0_140_2), .A4 (n_0_140_1));
NAND3_X1 i_0_123_31 (.ZN (n_0_123_30), .A1 (n_0_123_27), .A2 (n_0_123_28), .A3 (n_0_123_29));
NOR2_X1 i_0_123_30 (.ZN (n_0_123_29), .A1 (n_0_123_13), .A2 (n_0_123_23));
NOR2_X1 i_0_123_29 (.ZN (n_0_123_28), .A1 (n_0_123_22), .A2 (n_0_123_21));
NOR2_X1 i_0_123_28 (.ZN (n_0_123_27), .A1 (n_0_123_17), .A2 (n_0_123_20));
NOR2_X1 i_0_123_27 (.ZN (n_0_123_26), .A1 (n_0_123_17), .A2 (n_0_123_13));
NOR2_X1 i_0_123_26 (.ZN (n_0_123_25), .A1 (n_0_123_20), .A2 (n_0_123_21));
NOR2_X1 i_0_123_25 (.ZN (n_0_123_24), .A1 (n_0_123_22), .A2 (n_0_123_23));
NAND3_X1 i_0_123_24 (.ZN (n_0_123_23), .A1 (n_0_123_4), .A2 (n_0_123_2), .A3 (n_0_123_6));
NAND3_X1 i_0_123_23 (.ZN (n_0_123_22), .A1 (n_0_123_1), .A2 (n_0_123_3), .A3 (n_0_123_5));
NAND3_X1 i_0_123_22 (.ZN (n_0_123_21), .A1 (n_0_123_10), .A2 (n_0_123_8), .A3 (n_0_123_12));
NAND3_X1 i_0_123_21 (.ZN (n_0_123_20), .A1 (n_0_123_7), .A2 (n_0_123_9), .A3 (n_0_123_11));
NAND2_X1 i_0_123_20 (.ZN (n_0_123_19), .A1 (n_0_123_30), .A2 (\mem[5][11] ));
INV_X1 i_0_123_19 (.ZN (n_0_123_18), .A (sps__n112));
NAND4_X1 i_0_123_18 (.ZN (n_0_123_17), .A1 (n_0_123_18), .A2 (sps__n3), .A3 (sps__n121), .A4 (sps__n99));
INV_X1 i_0_123_17 (.ZN (n_0_123_16), .A (sps__n21));
INV_X1 i_0_123_16 (.ZN (n_0_123_15), .A (sps__n80));
INV_X1 i_0_123_15 (.ZN (n_0_123_14), .A (sps__n103));
NAND3_X1 i_0_123_14 (.ZN (n_0_123_13), .A1 (n_0_123_16), .A2 (n_0_123_15), .A3 (n_0_123_14));
INV_X1 i_0_123_13 (.ZN (n_0_123_12), .A (sps__n63));
INV_X1 i_0_123_12 (.ZN (n_0_123_11), .A (sps__n74));
INV_X1 i_0_123_11 (.ZN (n_0_123_10), .A (sps__n8));
INV_X1 i_0_123_10 (.ZN (n_0_123_9), .A (sps__n14));
INV_X1 i_0_123_9 (.ZN (n_0_123_8), .A (sps__n87));
INV_X1 i_0_123_8 (.ZN (n_0_123_7), .A (sps__n34));
INV_X1 i_0_123_7 (.ZN (n_0_123_6), .A (sps__n91));
INV_X1 i_0_123_6 (.ZN (n_0_123_5), .A (sps__n68));
INV_X1 i_0_123_5 (.ZN (n_0_123_4), .A (sps__n26));
INV_X1 i_0_123_4 (.ZN (n_0_123_3), .A (sps__n44));
INV_X1 i_0_123_3 (.ZN (n_0_123_2), .A (sps__n49));
INV_X1 i_0_123_2 (.ZN (n_0_123_1), .A (sps__n57));
NAND4_X1 i_0_123_1 (.ZN (n_0_123_0), .A1 (n_0_123_26), .A2 (n_0_123_25), .A3 (n_0_123_24), .A4 (data[11]));
NAND2_X1 i_0_123_0 (.ZN (n_0_80), .A1 (n_0_123_19), .A2 (n_0_123_0));
NAND3_X1 i_0_106_31 (.ZN (n_0_106_30), .A1 (n_0_106_27), .A2 (n_0_106_28), .A3 (n_0_106_29));
NOR2_X1 i_0_106_30 (.ZN (n_0_106_29), .A1 (n_0_106_13), .A2 (n_0_106_23));
NOR2_X1 i_0_106_29 (.ZN (n_0_106_28), .A1 (n_0_106_22), .A2 (n_0_106_21));
NOR2_X1 i_0_106_28 (.ZN (n_0_106_27), .A1 (n_0_106_17), .A2 (n_0_106_20));
NOR2_X1 i_0_106_27 (.ZN (n_0_106_26), .A1 (n_0_106_17), .A2 (n_0_106_13));
NOR2_X1 i_0_106_26 (.ZN (n_0_106_25), .A1 (n_0_106_20), .A2 (n_0_106_21));
NOR2_X1 i_0_106_25 (.ZN (n_0_106_24), .A1 (n_0_106_22), .A2 (n_0_106_23));
NAND3_X1 i_0_106_24 (.ZN (n_0_106_23), .A1 (n_0_106_4), .A2 (n_0_106_2), .A3 (n_0_106_6));
NAND3_X1 i_0_106_23 (.ZN (n_0_106_22), .A1 (n_0_106_1), .A2 (n_0_106_3), .A3 (n_0_106_5));
NAND3_X1 i_0_106_22 (.ZN (n_0_106_21), .A1 (n_0_106_10), .A2 (n_0_106_8), .A3 (n_0_106_12));
NAND3_X1 i_0_106_21 (.ZN (n_0_106_20), .A1 (n_0_106_7), .A2 (n_0_106_9), .A3 (n_0_106_11));
NAND2_X1 i_0_106_20 (.ZN (n_0_106_19), .A1 (n_0_106_30), .A2 (\mem[6][11] ));
INV_X1 i_0_106_19 (.ZN (n_0_106_18), .A (sps__n99));
NAND4_X1 i_0_106_18 (.ZN (n_0_106_17), .A1 (n_0_106_18), .A2 (sps__n3), .A3 (sps__n121), .A4 (sps__n112));
INV_X1 i_0_106_17 (.ZN (n_0_106_16), .A (sps__n19));
INV_X1 i_0_106_16 (.ZN (n_0_106_15), .A (sps__n81));
INV_X1 i_0_106_15 (.ZN (n_0_106_14), .A (sps__n104));
NAND3_X1 i_0_106_14 (.ZN (n_0_106_13), .A1 (n_0_106_16), .A2 (n_0_106_15), .A3 (n_0_106_14));
INV_X1 i_0_106_13 (.ZN (n_0_106_12), .A (sps__n62));
INV_X1 i_0_106_12 (.ZN (n_0_106_11), .A (sps__n74));
INV_X1 i_0_106_11 (.ZN (n_0_106_10), .A (sps__n8));
INV_X1 i_0_106_10 (.ZN (n_0_106_9), .A (sps__n14));
INV_X1 i_0_106_9 (.ZN (n_0_106_8), .A (sps__n86));
INV_X1 i_0_106_8 (.ZN (n_0_106_7), .A (sps__n34));
INV_X1 i_0_106_7 (.ZN (n_0_106_6), .A (sps__n91));
INV_X1 i_0_106_6 (.ZN (n_0_106_5), .A (sps__n68));
INV_X1 i_0_106_5 (.ZN (n_0_106_4), .A (sps__n28));
INV_X1 i_0_106_4 (.ZN (n_0_106_3), .A (sps__n44));
INV_X1 i_0_106_3 (.ZN (n_0_106_2), .A (sps__n50));
INV_X1 i_0_106_2 (.ZN (n_0_106_1), .A (sps__n55));
NAND4_X1 i_0_106_1 (.ZN (n_0_106_0), .A1 (n_0_106_26), .A2 (n_0_106_25), .A3 (n_0_106_24), .A4 (data[11]));
NAND2_X1 i_0_106_0 (.ZN (n_0_79), .A1 (n_0_106_19), .A2 (n_0_106_0));
NAND3_X1 i_0_89_27 (.ZN (n_0_89_26), .A1 (n_0_89_23), .A2 (n_0_89_24), .A3 (n_0_89_25));
NOR2_X1 i_0_89_26 (.ZN (n_0_89_25), .A1 (n_0_89_17), .A2 (n_0_89_13));
NOR2_X1 i_0_89_25 (.ZN (n_0_89_24), .A1 (n_0_89_19), .A2 (n_0_89_20));
NOR2_X1 i_0_89_24 (.ZN (n_0_89_23), .A1 (n_0_89_21), .A2 (n_0_89_22));
NAND3_X1 i_0_89_23 (.ZN (n_0_89_22), .A1 (n_0_89_4), .A2 (n_0_89_2), .A3 (n_0_89_6));
NAND3_X1 i_0_89_22 (.ZN (n_0_89_21), .A1 (n_0_89_1), .A2 (n_0_89_3), .A3 (n_0_89_5));
NAND3_X1 i_0_89_21 (.ZN (n_0_89_20), .A1 (n_0_89_10), .A2 (n_0_89_8), .A3 (n_0_89_12));
NAND3_X1 i_0_89_20 (.ZN (n_0_89_19), .A1 (n_0_89_7), .A2 (n_0_89_9), .A3 (n_0_89_11));
NAND2_X1 i_0_89_19 (.ZN (n_0_89_18), .A1 (n_0_89_26), .A2 (\mem[7][11] ));
NAND4_X1 i_0_89_18 (.ZN (n_0_89_17), .A1 (sps__n2), .A2 (sps__n121), .A3 (sps__n114), .A4 (sps__n97));
INV_X1 i_0_89_17 (.ZN (n_0_89_16), .A (sps__n20));
INV_X1 i_0_89_16 (.ZN (n_0_89_15), .A (sps__n80));
INV_X1 i_0_89_15 (.ZN (n_0_89_14), .A (sps__n103));
NAND3_X1 i_0_89_14 (.ZN (n_0_89_13), .A1 (n_0_89_16), .A2 (n_0_89_15), .A3 (n_0_89_14));
INV_X1 i_0_89_13 (.ZN (n_0_89_12), .A (sps__n61));
INV_X1 i_0_89_12 (.ZN (n_0_89_11), .A (sps__n74));
INV_X1 i_0_89_11 (.ZN (n_0_89_10), .A (sps__n8));
INV_X1 i_0_89_10 (.ZN (n_0_89_9), .A (sps__n14));
INV_X1 i_0_89_9 (.ZN (n_0_89_8), .A (sps__n85));
INV_X1 i_0_89_8 (.ZN (n_0_89_7), .A (sps__n36));
INV_X1 i_0_89_7 (.ZN (n_0_89_6), .A (sps__n91));
INV_X1 i_0_89_6 (.ZN (n_0_89_5), .A (sps__n68));
INV_X1 i_0_89_5 (.ZN (n_0_89_4), .A (sps__n26));
INV_X1 i_0_89_4 (.ZN (n_0_89_3), .A (sps__n44));
INV_X1 i_0_89_3 (.ZN (n_0_89_2), .A (sps__n50));
INV_X1 i_0_89_2 (.ZN (n_0_89_1), .A (sps__n55));
NAND4_X1 i_0_89_1 (.ZN (n_0_89_0), .A1 (n_0_89_25), .A2 (n_0_89_24), .A3 (n_0_89_23), .A4 (data[11]));
NAND2_X1 i_0_89_0 (.ZN (n_0_78), .A1 (n_0_89_18), .A2 (n_0_89_0));
NAND3_X1 i_0_72_35 (.ZN (n_0_77), .A1 (n_0_72_32), .A2 (n_0_72_33), .A3 (n_0_72_34));
NAND2_X1 i_0_72_34 (.ZN (n_0_72_34), .A1 (n_0_72_23), .A2 (\mem[8][11] ));
NAND3_X1 i_0_72_29 (.ZN (n_0_72_33), .A1 (n_0_72_26), .A2 (n_0_72_31), .A3 (n_0_72_28));
NAND2_X1 i_0_72_28 (.ZN (n_0_72_32), .A1 (n_0_72_27), .A2 (\mem[8][11] ));
NOR2_X1 i_0_72_24 (.ZN (n_0_72_31), .A1 (n_0_72_18), .A2 (n_0_72_0));
INV_X1 i_0_72_23 (.ZN (n_0_72_30), .A (n_0_72_0));
INV_X1 i_0_72_22 (.ZN (n_0_72_29), .A (n_0_72_18));
INV_X1 i_0_72_21 (.ZN (n_0_72_28), .A (n_0_72_5));
NAND3_X1 i_0_72_20 (.ZN (n_0_72_27), .A1 (n_0_72_28), .A2 (n_0_72_30), .A3 (n_0_72_9));
NOR2_X1 i_0_72_19 (.ZN (n_0_72_26), .A1 (n_0_72_14), .A2 (n_0_72_24));
INV_X1 i_0_72_18 (.ZN (n_0_72_25), .A (n_0_72_14));
NAND2_X1 i_0_72_17 (.ZN (n_0_72_24), .A1 (n_0_72_9), .A2 (data[11]));
NAND2_X1 i_0_72_16 (.ZN (n_0_72_23), .A1 (n_0_72_29), .A2 (n_0_72_25));
INV_X1 i_0_72_33 (.ZN (n_0_72_22), .A (sps__n36));
INV_X1 i_0_72_32 (.ZN (n_0_72_21), .A (sps__n8));
INV_X1 i_0_72_31 (.ZN (n_0_72_20), .A (sps__n14));
INV_X1 i_0_72_30 (.ZN (n_0_72_19), .A (sps__n50));
NAND4_X1 i_0_72_3 (.ZN (n_0_72_18), .A1 (n_0_72_22), .A2 (n_0_72_21), .A3 (n_0_72_20), .A4 (n_0_72_19));
INV_X1 i_0_72_27 (.ZN (n_0_72_17), .A (sps__n62));
INV_X1 i_0_72_26 (.ZN (n_0_72_16), .A (sps__n74));
INV_X1 i_0_72_25 (.ZN (n_0_72_15), .A (sps__n86));
NAND4_X1 i_0_72_8 (.ZN (n_0_72_14), .A1 (n_0_72_17), .A2 (n_0_72_16), .A3 (n_0_72_15), .A4 (sps__n2));
INV_X1 i_0_72_15 (.ZN (n_0_72_13), .A (sps__n121));
INV_X1 i_0_72_14 (.ZN (n_0_72_12), .A (sps__n114));
INV_X1 i_0_72_13 (.ZN (n_0_72_11), .A (sps__n97));
NAND3_X1 i_0_72_12 (.ZN (n_0_72_10), .A1 (n_0_72_13), .A2 (n_0_72_12), .A3 (n_0_72_11));
INV_X1 i_0_72_11 (.ZN (n_0_72_9), .A (n_0_72_10));
INV_X1 i_0_72_10 (.ZN (n_0_72_8), .A (sps__n68));
INV_X1 i_0_72_9 (.ZN (n_0_72_7), .A (sps__n20));
INV_X1 i_0_72_7 (.ZN (n_0_72_6), .A (sps__n80));
NAND4_X1 i_0_72_6 (.ZN (n_0_72_5), .A1 (n_0_72_8), .A2 (n_0_72_7), .A3 (n_0_72_6), .A4 (sps__n104));
INV_X1 i_0_72_5 (.ZN (n_0_72_4), .A (sps__n55));
INV_X1 i_0_72_4 (.ZN (n_0_72_3), .A (sps__n26));
INV_X1 i_0_72_2 (.ZN (n_0_72_2), .A (sps__n44));
INV_X1 i_0_72_1 (.ZN (n_0_72_1), .A (sps__n91));
NAND4_X1 i_0_72_0 (.ZN (n_0_72_0), .A1 (n_0_72_4), .A2 (n_0_72_3), .A3 (n_0_72_2), .A4 (n_0_72_1));
NOR2_X1 i_0_55_34 (.ZN (n_0_55_33), .A1 (n_0_55_19), .A2 (n_0_55_0));
INV_X1 i_0_55_33 (.ZN (n_0_55_32), .A (n_0_55_0));
INV_X1 i_0_55_28 (.ZN (n_0_55_31), .A (n_0_55_19));
NAND2_X1 i_0_55_27 (.ZN (n_0_55_30), .A1 (n_0_55_29), .A2 (\mem[9][11] ));
NAND3_X1 i_0_55_23 (.ZN (n_0_55_29), .A1 (n_0_55_5), .A2 (n_0_55_32), .A3 (n_0_55_10));
NAND3_X1 i_0_55_22 (.ZN (n_0_55_28), .A1 (n_0_55_27), .A2 (n_0_55_33), .A3 (n_0_55_14));
NOR2_X1 i_0_55_21 (.ZN (n_0_55_27), .A1 (n_0_55_6), .A2 (n_0_55_26));
NAND2_X1 i_0_55_20 (.ZN (n_0_55_26), .A1 (n_0_55_10), .A2 (data[11]));
NAND2_X1 i_0_55_19 (.ZN (n_0_55_25), .A1 (n_0_55_31), .A2 (n_0_55_14));
NAND3_X1 i_0_55_18 (.ZN (n_0_76), .A1 (n_0_55_28), .A2 (n_0_55_30), .A3 (n_0_55_24));
NAND2_X1 i_0_55_17 (.ZN (n_0_55_24), .A1 (n_0_55_25), .A2 (\mem[9][11] ));
INV_X1 i_0_55_32 (.ZN (n_0_55_23), .A (sps__n35));
INV_X1 i_0_55_31 (.ZN (n_0_55_22), .A (sps__n8));
INV_X1 i_0_55_30 (.ZN (n_0_55_21), .A (sps__n13));
INV_X1 i_0_55_29 (.ZN (n_0_55_20), .A (sps__n49));
NAND4_X1 i_0_55_3 (.ZN (n_0_55_19), .A1 (n_0_55_23), .A2 (n_0_55_22), .A3 (n_0_55_21), .A4 (n_0_55_20));
INV_X1 i_0_55_26 (.ZN (n_0_55_18), .A (sps__n63));
INV_X1 i_0_55_25 (.ZN (n_0_55_17), .A (sps__n74));
INV_X1 i_0_55_24 (.ZN (n_0_55_16), .A (sps__n87));
NAND4_X1 i_0_55_6 (.ZN (n_0_55_15), .A1 (n_0_55_18), .A2 (n_0_55_17), .A3 (n_0_55_16), .A4 (sps__n1));
INV_X1 i_0_55_16 (.ZN (n_0_55_14), .A (n_0_55_15));
INV_X1 i_0_55_15 (.ZN (n_0_55_13), .A (sps__n121));
INV_X1 i_0_55_14 (.ZN (n_0_55_12), .A (sps__n112));
NAND3_X1 i_0_55_13 (.ZN (n_0_55_11), .A1 (n_0_55_13), .A2 (n_0_55_12), .A3 (sps__n97));
INV_X1 i_0_55_12 (.ZN (n_0_55_10), .A (n_0_55_11));
INV_X1 i_0_55_11 (.ZN (n_0_55_9), .A (sps__n68));
INV_X1 i_0_55_10 (.ZN (n_0_55_8), .A (sps__n21));
INV_X1 i_0_55_9 (.ZN (n_0_55_7), .A (sps__n80));
NAND4_X1 i_0_55_8 (.ZN (n_0_55_6), .A1 (n_0_55_9), .A2 (n_0_55_8), .A3 (n_0_55_7), .A4 (sps__n103));
INV_X1 i_0_55_7 (.ZN (n_0_55_5), .A (n_0_55_6));
INV_X1 i_0_55_5 (.ZN (n_0_55_4), .A (sps__n57));
INV_X1 i_0_55_4 (.ZN (n_0_55_3), .A (sps__n27));
INV_X1 i_0_55_2 (.ZN (n_0_55_2), .A (sps__n44));
INV_X1 i_0_55_1 (.ZN (n_0_55_1), .A (sps__n93));
NAND4_X1 i_0_55_0 (.ZN (n_0_55_0), .A1 (n_0_55_4), .A2 (n_0_55_3), .A3 (n_0_55_2), .A4 (n_0_55_1));
NOR2_X1 i_0_38_34 (.ZN (n_0_38_33), .A1 (n_0_38_19), .A2 (n_0_38_0));
INV_X1 i_0_38_33 (.ZN (n_0_38_32), .A (n_0_38_0));
INV_X1 i_0_38_28 (.ZN (n_0_38_31), .A (n_0_38_19));
NAND2_X1 i_0_38_27 (.ZN (n_0_38_30), .A1 (n_0_38_29), .A2 (\mem[10][11] ));
NAND3_X1 i_0_38_23 (.ZN (n_0_38_29), .A1 (n_0_38_5), .A2 (n_0_38_32), .A3 (n_0_38_10));
NAND3_X1 i_0_38_22 (.ZN (n_0_38_28), .A1 (n_0_38_27), .A2 (n_0_38_33), .A3 (n_0_38_14));
NOR2_X1 i_0_38_21 (.ZN (n_0_38_27), .A1 (n_0_38_6), .A2 (n_0_38_26));
NAND2_X1 i_0_38_20 (.ZN (n_0_38_26), .A1 (n_0_38_10), .A2 (data[11]));
NAND2_X1 i_0_38_19 (.ZN (n_0_38_25), .A1 (n_0_38_31), .A2 (n_0_38_14));
NAND3_X1 i_0_38_18 (.ZN (n_0_75), .A1 (n_0_38_28), .A2 (n_0_38_30), .A3 (n_0_38_24));
NAND2_X1 i_0_38_17 (.ZN (n_0_38_24), .A1 (n_0_38_25), .A2 (\mem[10][11] ));
INV_X1 i_0_38_32 (.ZN (n_0_38_23), .A (sps__n36));
INV_X1 i_0_38_31 (.ZN (n_0_38_22), .A (sps__n8));
INV_X1 i_0_38_30 (.ZN (n_0_38_21), .A (sps__n14));
INV_X1 i_0_38_29 (.ZN (n_0_38_20), .A (sps__n50));
NAND4_X1 i_0_38_3 (.ZN (n_0_38_19), .A1 (n_0_38_23), .A2 (n_0_38_22), .A3 (n_0_38_21), .A4 (n_0_38_20));
INV_X1 i_0_38_26 (.ZN (n_0_38_18), .A (sps__n62));
INV_X1 i_0_38_25 (.ZN (n_0_38_17), .A (sps__n74));
INV_X1 i_0_38_24 (.ZN (n_0_38_16), .A (sps__n85));
NAND4_X1 i_0_38_6 (.ZN (n_0_38_15), .A1 (n_0_38_18), .A2 (n_0_38_17), .A3 (n_0_38_16), .A4 (sps__n2));
INV_X1 i_0_38_16 (.ZN (n_0_38_14), .A (n_0_38_15));
INV_X1 i_0_38_15 (.ZN (n_0_38_13), .A (sps__n121));
INV_X1 i_0_38_14 (.ZN (n_0_38_12), .A (sps__n97));
NAND3_X1 i_0_38_13 (.ZN (n_0_38_11), .A1 (n_0_38_13), .A2 (n_0_38_12), .A3 (sps__n114));
INV_X1 i_0_38_12 (.ZN (n_0_38_10), .A (n_0_38_11));
INV_X1 i_0_38_11 (.ZN (n_0_38_9), .A (sps__n68));
INV_X1 i_0_38_10 (.ZN (n_0_38_8), .A (sps__n20));
INV_X1 i_0_38_9 (.ZN (n_0_38_7), .A (sps__n81));
NAND4_X1 i_0_38_8 (.ZN (n_0_38_6), .A1 (n_0_38_9), .A2 (n_0_38_8), .A3 (n_0_38_7), .A4 (sps__n104));
INV_X1 i_0_38_7 (.ZN (n_0_38_5), .A (n_0_38_6));
INV_X1 i_0_38_5 (.ZN (n_0_38_4), .A (sps__n55));
INV_X1 i_0_38_4 (.ZN (n_0_38_3), .A (sps__n26));
INV_X1 i_0_38_2 (.ZN (n_0_38_2), .A (sps__n44));
INV_X1 i_0_38_1 (.ZN (n_0_38_1), .A (sps__n91));
NAND4_X1 i_0_38_0 (.ZN (n_0_38_0), .A1 (n_0_38_4), .A2 (n_0_38_3), .A3 (n_0_38_2), .A4 (n_0_38_1));
INV_X1 i_0_21_37 (.ZN (n_0_21_36), .A (sps__n114));
INV_X1 i_0_21_36 (.ZN (n_0_21_35), .A (sps__n103));
NAND3_X1 i_0_21_35 (.ZN (n_0_21_34), .A1 (n_0_21_35), .A2 (\mem[5][12] ), .A3 (sps__n123));
INV_X1 i_0_21_34 (.ZN (n_0_21_33), .A (sps__n123));
INV_X1 i_0_21_33 (.ZN (n_0_21_32), .A (\mem[1][12] ));
NAND2_X1 i_0_21_32 (.ZN (n_0_21_31), .A1 (n_0_21_35), .A2 (n_0_21_32));
INV_X1 i_0_21_31 (.ZN (n_0_21_30), .A (\mem[9][12] ));
NAND2_X1 i_0_21_30 (.ZN (n_0_21_29), .A1 (sps__n103), .A2 (n_0_21_30));
NAND3_X1 i_0_21_29 (.ZN (n_0_21_28), .A1 (n_0_21_31), .A2 (n_0_21_33), .A3 (n_0_21_29));
NAND3_X1 i_0_21_28 (.ZN (n_0_21_27), .A1 (n_0_21_28), .A2 (n_0_21_36), .A3 (n_0_21_34));
INV_X1 i_0_21_27 (.ZN (n_0_21_26), .A (\mem[3][12] ));
NAND2_X1 i_0_21_26 (.ZN (n_0_21_25), .A1 (n_0_21_33), .A2 (n_0_21_26));
INV_X1 i_0_21_24 (.ZN (n_0_21_24), .A (\mem[7][12] ));
NAND2_X1 i_0_21_23 (.ZN (n_0_21_23), .A1 (sps__n123), .A2 (n_0_21_24));
NAND3_X1 i_0_21_22 (.ZN (n_0_21_22), .A1 (n_0_21_25), .A2 (n_0_21_35), .A3 (n_0_21_23));
NAND2_X1 i_0_21_21 (.ZN (n_0_21_21), .A1 (n_0_21_22), .A2 (sps__n114));
NAND3_X1 i_0_21_20 (.ZN (n_0_21_19), .A1 (n_0_21_27), .A2 (sps__n98), .A3 (n_0_21_21));
INV_X1 i_0_21_19 (.ZN (n_0_21_18), .A (sps__n98));
INV_X1 i_0_21_18 (.ZN (n_0_21_17), .A (\mem[8][12] ));
NAND2_X1 i_0_21_17 (.ZN (n_0_21_16), .A1 (n_0_21_36), .A2 (n_0_21_17));
INV_X1 i_0_21_16 (.ZN (n_0_21_15), .A (\mem[10][12] ));
NAND2_X1 i_0_21_15 (.ZN (n_0_21_14), .A1 (sps__n114), .A2 (n_0_21_15));
NAND3_X1 i_0_21_14 (.ZN (n_0_21_13), .A1 (n_0_21_16), .A2 (n_0_21_33), .A3 (n_0_21_14));
NAND2_X1 i_0_21_13 (.ZN (n_0_21_12), .A1 (n_0_21_13), .A2 (sps__n103));
NAND2_X1 i_0_21_12 (.ZN (n_0_21_11), .A1 (n_0_21_36), .A2 (\mem[0][12] ));
NAND2_X1 i_0_21_11 (.ZN (n_0_21_10), .A1 (sps__n114), .A2 (\mem[2][12] ));
NAND4_X1 i_0_21_10 (.ZN (n_0_21_9), .A1 (n_0_21_11), .A2 (n_0_21_10), .A3 (n_0_21_35), .A4 (n_0_21_33));
NAND2_X1 i_0_21_9 (.ZN (n_0_21_8), .A1 (n_0_21_36), .A2 (\mem[4][12] ));
NAND2_X1 i_0_21_8 (.ZN (n_0_21_7), .A1 (sps__n114), .A2 (\mem[6][12] ));
NAND3_X1 i_0_21_7 (.ZN (n_0_21_6), .A1 (n_0_21_8), .A2 (sps__n123), .A3 (n_0_21_7));
NAND4_X1 i_0_21_6 (.ZN (n_0_21_5), .A1 (n_0_21_12), .A2 (n_0_21_18), .A3 (n_0_21_9), .A4 (n_0_21_6));
NAND2_X1 i_0_21_5 (.ZN (n_0_21_4), .A1 (n_0_21_5), .A2 (n_0_21_19));
NAND2_X1 i_0_21_4 (.ZN (n_0_21_3), .A1 (n_0_21_4), .A2 (n_0_5));
INV_X1 i_0_21_3 (.ZN (n_0_21_2), .A (n_0_5));
INV_X1 i_0_21_2 (.ZN (n_0_21_1), .A (n_0_21_20));
NAND2_X1 i_0_21_1 (.ZN (n_0_21_0), .A1 (n_0_21_2), .A2 (n_0_21_1));
NAND2_X1 i_0_21_0 (.ZN (n_0_71), .A1 (n_0_21_0), .A2 (n_0_21_3));
INV_X1 i_0_21_25 (.ZN (n_0_21_20), .A (dataout[12]));
NAND3_X1 i_0_3_37 (.ZN (n_0_64), .A1 (n_0_3_34), .A2 (n_0_3_35), .A3 (n_0_3_36));
NAND2_X1 i_0_3_36 (.ZN (n_0_3_36), .A1 (n_0_3_25), .A2 (\mem[0][12] ));
NAND3_X1 i_0_3_35 (.ZN (n_0_3_35), .A1 (n_0_3_27), .A2 (n_0_3_33), .A3 (n_0_3_30));
NAND2_X1 i_0_3_34 (.ZN (n_0_3_34), .A1 (n_0_3_24), .A2 (\mem[0][12] ));
NOR2_X1 i_0_3_33 (.ZN (n_0_3_33), .A1 (n_0_3_0), .A2 (n_0_3_19));
INV_X1 i_0_3_32 (.ZN (n_0_3_32), .A (n_0_3_19));
INV_X1 i_0_3_31 (.ZN (n_0_3_31), .A (n_0_3_0));
NOR2_X1 i_0_3_30 (.ZN (n_0_3_30), .A1 (n_0_3_5), .A2 (n_0_3_15));
INV_X1 i_0_3_29 (.ZN (n_0_3_29), .A (n_0_3_15));
INV_X1 i_0_3_28 (.ZN (n_0_3_28), .A (n_0_3_5));
INV_X1 i_0_3_27 (.ZN (n_0_3_27), .A (n_0_3_26));
NAND2_X1 i_0_3_26 (.ZN (n_0_3_26), .A1 (n_0_3_10), .A2 (data[12]));
NAND2_X1 i_0_3_25 (.ZN (n_0_3_25), .A1 (n_0_3_31), .A2 (n_0_3_28));
NAND3_X1 i_0_3_24 (.ZN (n_0_3_24), .A1 (n_0_3_32), .A2 (n_0_3_29), .A3 (n_0_3_10));
INV_X1 i_0_3_23 (.ZN (n_0_3_23), .A (sps__n36));
INV_X1 i_0_3_22 (.ZN (n_0_3_22), .A (sps__n7));
INV_X1 i_0_3_21 (.ZN (n_0_3_21), .A (sps__n14));
INV_X1 i_0_3_20 (.ZN (n_0_3_20), .A (sps__n51));
NAND4_X1 i_0_3_19 (.ZN (n_0_3_19), .A1 (n_0_3_23), .A2 (n_0_3_22), .A3 (n_0_3_21), .A4 (n_0_3_20));
INV_X1 i_0_3_18 (.ZN (n_0_3_18), .A (sps__n62));
INV_X1 i_0_3_17 (.ZN (n_0_3_17), .A (sps__n74));
INV_X1 i_0_3_12 (.ZN (n_0_3_16), .A (sps__n86));
NAND4_X1 i_0_3_11 (.ZN (n_0_3_15), .A1 (n_0_3_18), .A2 (n_0_3_17), .A3 (n_0_3_16), .A4 (sps__n2));
INV_X1 i_0_3_6 (.ZN (n_0_3_14), .A (sps__n123));
INV_X1 i_0_3_5 (.ZN (n_0_3_13), .A (sps__n114));
INV_X1 i_0_3_4 (.ZN (n_0_3_12), .A (sps__n98));
NAND3_X1 i_0_3_1 (.ZN (n_0_3_11), .A1 (n_0_3_14), .A2 (n_0_3_13), .A3 (n_0_3_12));
INV_X1 i_0_3_0 (.ZN (n_0_3_10), .A (n_0_3_11));
INV_X1 i_0_3_16 (.ZN (n_0_3_9), .A (sps__n68));
INV_X1 i_0_3_15 (.ZN (n_0_3_8), .A (sps__n20));
INV_X1 i_0_3_14 (.ZN (n_0_3_7), .A (sps__n80));
INV_X1 i_0_3_13 (.ZN (n_0_3_6), .A (sps__n103));
NAND4_X1 i_0_3_3 (.ZN (n_0_3_5), .A1 (n_0_3_9), .A2 (n_0_3_8), .A3 (n_0_3_7), .A4 (n_0_3_6));
INV_X1 i_0_3_10 (.ZN (n_0_3_4), .A (sps__n55));
INV_X1 i_0_3_9 (.ZN (n_0_3_3), .A (address[9]));
INV_X1 i_0_3_8 (.ZN (n_0_3_2), .A (sps__n42));
INV_X1 i_0_3_7 (.ZN (n_0_3_1), .A (sps__n92));
NAND4_X1 i_0_3_2 (.ZN (n_0_3_0), .A1 (n_0_3_4), .A2 (n_0_3_3), .A3 (n_0_3_2), .A4 (n_0_3_1));
NAND3_X1 i_0_67_36 (.ZN (n_0_63), .A1 (n_0_67_33), .A2 (n_0_67_34), .A3 (n_0_67_35));
NAND2_X1 i_0_67_35 (.ZN (n_0_67_35), .A1 (n_0_67_24), .A2 (\mem[1][12] ));
NAND2_X1 i_0_67_34 (.ZN (n_0_67_34), .A1 (n_0_67_23), .A2 (\mem[1][12] ));
NAND3_X1 i_0_67_33 (.ZN (n_0_67_33), .A1 (n_0_67_26), .A2 (n_0_67_32), .A3 (n_0_67_29));
NOR2_X1 i_0_67_32 (.ZN (n_0_67_32), .A1 (n_0_67_0), .A2 (n_0_67_18));
INV_X1 i_0_67_31 (.ZN (n_0_67_31), .A (n_0_67_18));
INV_X1 i_0_67_30 (.ZN (n_0_67_30), .A (n_0_67_0));
NOR2_X1 i_0_67_29 (.ZN (n_0_67_29), .A1 (n_0_67_5), .A2 (n_0_67_14));
INV_X1 i_0_67_28 (.ZN (n_0_67_28), .A (n_0_67_14));
INV_X1 i_0_67_27 (.ZN (n_0_67_27), .A (n_0_67_5));
INV_X1 i_0_67_26 (.ZN (n_0_67_26), .A (n_0_67_25));
NAND2_X1 i_0_67_25 (.ZN (n_0_67_25), .A1 (n_0_67_10), .A2 (data[12]));
NAND2_X1 i_0_67_24 (.ZN (n_0_67_24), .A1 (n_0_67_30), .A2 (n_0_67_27));
NAND3_X1 i_0_67_23 (.ZN (n_0_67_23), .A1 (n_0_67_31), .A2 (n_0_67_28), .A3 (n_0_67_10));
INV_X1 i_0_67_22 (.ZN (n_0_67_22), .A (sps__n36));
INV_X1 i_0_67_21 (.ZN (n_0_67_21), .A (sps__n7));
INV_X1 i_0_67_20 (.ZN (n_0_67_20), .A (sps__n14));
INV_X1 i_0_67_19 (.ZN (n_0_67_19), .A (sps__n50));
NAND4_X1 i_0_67_18 (.ZN (n_0_67_18), .A1 (n_0_67_22), .A2 (n_0_67_21), .A3 (n_0_67_20), .A4 (n_0_67_19));
INV_X1 i_0_67_17 (.ZN (n_0_67_17), .A (sps__n62));
INV_X1 i_0_67_12 (.ZN (n_0_67_16), .A (sps__n74));
INV_X1 i_0_67_11 (.ZN (n_0_67_15), .A (sps__n86));
NAND4_X1 i_0_67_6 (.ZN (n_0_67_14), .A1 (n_0_67_17), .A2 (n_0_67_16), .A3 (n_0_67_15), .A4 (sps__n2));
INV_X1 i_0_67_5 (.ZN (n_0_67_13), .A (sps__n123));
INV_X1 i_0_67_4 (.ZN (n_0_67_12), .A (sps__n114));
NAND3_X1 i_0_67_1 (.ZN (n_0_67_11), .A1 (n_0_67_13), .A2 (n_0_67_12), .A3 (sps__n98));
INV_X1 i_0_67_0 (.ZN (n_0_67_10), .A (n_0_67_11));
INV_X1 i_0_67_16 (.ZN (n_0_67_9), .A (sps__n69));
INV_X1 i_0_67_15 (.ZN (n_0_67_8), .A (sps__n20));
INV_X1 i_0_67_14 (.ZN (n_0_67_7), .A (address[4]));
INV_X1 i_0_67_13 (.ZN (n_0_67_6), .A (sps__n103));
NAND4_X1 i_0_67_3 (.ZN (n_0_67_5), .A1 (n_0_67_9), .A2 (n_0_67_8), .A3 (n_0_67_7), .A4 (n_0_67_6));
INV_X1 i_0_67_10 (.ZN (n_0_67_4), .A (sps__n55));
INV_X1 i_0_67_9 (.ZN (n_0_67_3), .A (address[9]));
INV_X1 i_0_67_8 (.ZN (n_0_67_2), .A (sps__n42));
INV_X1 i_0_67_7 (.ZN (n_0_67_1), .A (sps__n92));
NAND4_X1 i_0_67_2 (.ZN (n_0_67_0), .A1 (n_0_67_4), .A2 (n_0_67_3), .A3 (n_0_67_2), .A4 (n_0_67_1));
NAND3_X1 i_0_173_36 (.ZN (n_0_62), .A1 (n_0_173_33), .A2 (n_0_173_34), .A3 (n_0_173_35));
NAND2_X1 i_0_173_35 (.ZN (n_0_173_35), .A1 (n_0_173_24), .A2 (\mem[2][12] ));
NAND2_X1 i_0_173_34 (.ZN (n_0_173_34), .A1 (n_0_173_23), .A2 (\mem[2][12] ));
NAND3_X1 i_0_173_33 (.ZN (n_0_173_33), .A1 (n_0_173_26), .A2 (n_0_173_32), .A3 (n_0_173_29));
NOR2_X1 i_0_173_32 (.ZN (n_0_173_32), .A1 (n_0_173_0), .A2 (n_0_173_18));
INV_X1 i_0_173_31 (.ZN (n_0_173_31), .A (n_0_173_18));
INV_X1 i_0_173_30 (.ZN (n_0_173_30), .A (n_0_173_0));
NOR2_X1 i_0_173_29 (.ZN (n_0_173_29), .A1 (n_0_173_5), .A2 (n_0_173_14));
INV_X1 i_0_173_28 (.ZN (n_0_173_28), .A (n_0_173_14));
INV_X1 i_0_173_27 (.ZN (n_0_173_27), .A (n_0_173_5));
INV_X1 i_0_173_26 (.ZN (n_0_173_26), .A (n_0_173_25));
NAND2_X1 i_0_173_25 (.ZN (n_0_173_25), .A1 (n_0_173_10), .A2 (data[12]));
NAND2_X1 i_0_173_24 (.ZN (n_0_173_24), .A1 (n_0_173_30), .A2 (n_0_173_27));
NAND3_X1 i_0_173_23 (.ZN (n_0_173_23), .A1 (n_0_173_31), .A2 (n_0_173_28), .A3 (n_0_173_10));
INV_X1 i_0_173_22 (.ZN (n_0_173_22), .A (sps__n36));
INV_X1 i_0_173_21 (.ZN (n_0_173_21), .A (sps__n7));
INV_X1 i_0_173_20 (.ZN (n_0_173_20), .A (sps__n14));
INV_X1 i_0_173_19 (.ZN (n_0_173_19), .A (sps__n50));
NAND4_X1 i_0_173_18 (.ZN (n_0_173_18), .A1 (n_0_173_22), .A2 (n_0_173_21), .A3 (n_0_173_20), .A4 (n_0_173_19));
INV_X1 i_0_173_17 (.ZN (n_0_173_17), .A (RST));
INV_X1 i_0_173_12 (.ZN (n_0_173_16), .A (sps__n74));
INV_X1 i_0_173_11 (.ZN (n_0_173_15), .A (sps__n85));
NAND4_X1 i_0_173_6 (.ZN (n_0_173_14), .A1 (n_0_173_17), .A2 (n_0_173_16), .A3 (n_0_173_15), .A4 (sps__n2));
INV_X1 i_0_173_5 (.ZN (n_0_173_13), .A (sps__n123));
INV_X1 i_0_173_4 (.ZN (n_0_173_12), .A (sps__n98));
NAND3_X1 i_0_173_1 (.ZN (n_0_173_11), .A1 (n_0_173_13), .A2 (n_0_173_12), .A3 (sps__n114));
INV_X1 i_0_173_0 (.ZN (n_0_173_10), .A (n_0_173_11));
INV_X1 i_0_173_16 (.ZN (n_0_173_9), .A (sps__n69));
INV_X1 i_0_173_15 (.ZN (n_0_173_8), .A (sps__n20));
INV_X1 i_0_173_14 (.ZN (n_0_173_7), .A (address[4]));
INV_X1 i_0_173_13 (.ZN (n_0_173_6), .A (sps__n103));
NAND4_X1 i_0_173_3 (.ZN (n_0_173_5), .A1 (n_0_173_9), .A2 (n_0_173_8), .A3 (n_0_173_7), .A4 (n_0_173_6));
INV_X1 i_0_173_10 (.ZN (n_0_173_4), .A (sps__n56));
INV_X1 i_0_173_9 (.ZN (n_0_173_3), .A (sps__n26));
INV_X1 i_0_173_8 (.ZN (n_0_173_2), .A (sps__n42));
INV_X1 i_0_173_7 (.ZN (n_0_173_1), .A (sps__n91));
NAND4_X1 i_0_173_2 (.ZN (n_0_173_0), .A1 (n_0_173_4), .A2 (n_0_173_3), .A3 (n_0_173_2), .A4 (n_0_173_1));
NAND3_X1 i_0_156_31 (.ZN (n_0_156_30), .A1 (n_0_156_27), .A2 (n_0_156_28), .A3 (n_0_156_29));
NOR2_X1 i_0_156_30 (.ZN (n_0_156_29), .A1 (n_0_156_13), .A2 (n_0_156_23));
NOR2_X1 i_0_156_29 (.ZN (n_0_156_28), .A1 (n_0_156_22), .A2 (n_0_156_21));
NOR2_X1 i_0_156_28 (.ZN (n_0_156_27), .A1 (n_0_156_17), .A2 (n_0_156_20));
NOR2_X1 i_0_156_27 (.ZN (n_0_156_26), .A1 (n_0_156_17), .A2 (n_0_156_13));
NOR2_X1 i_0_156_26 (.ZN (n_0_156_25), .A1 (n_0_156_20), .A2 (n_0_156_21));
NOR2_X1 i_0_156_25 (.ZN (n_0_156_24), .A1 (n_0_156_22), .A2 (n_0_156_23));
NAND3_X1 i_0_156_24 (.ZN (n_0_156_23), .A1 (n_0_156_4), .A2 (n_0_156_2), .A3 (n_0_156_6));
NAND3_X1 i_0_156_23 (.ZN (n_0_156_22), .A1 (n_0_156_1), .A2 (n_0_156_3), .A3 (n_0_156_5));
NAND3_X1 i_0_156_22 (.ZN (n_0_156_21), .A1 (n_0_156_10), .A2 (n_0_156_8), .A3 (n_0_156_12));
NAND3_X1 i_0_156_21 (.ZN (n_0_156_20), .A1 (n_0_156_7), .A2 (n_0_156_9), .A3 (n_0_156_11));
NAND2_X1 i_0_156_20 (.ZN (n_0_156_19), .A1 (n_0_156_30), .A2 (\mem[3][12] ));
INV_X1 i_0_156_19 (.ZN (n_0_156_18), .A (sps__n123));
NAND4_X1 i_0_156_18 (.ZN (n_0_156_17), .A1 (n_0_156_18), .A2 (sps__n2), .A3 (sps__n114), .A4 (sps__n98));
INV_X1 i_0_156_17 (.ZN (n_0_156_16), .A (sps__n20));
INV_X1 i_0_156_16 (.ZN (n_0_156_15), .A (address[4]));
INV_X1 i_0_156_15 (.ZN (n_0_156_14), .A (sps__n103));
NAND3_X1 i_0_156_14 (.ZN (n_0_156_13), .A1 (n_0_156_16), .A2 (n_0_156_15), .A3 (n_0_156_14));
INV_X1 i_0_156_13 (.ZN (n_0_156_12), .A (RST));
INV_X1 i_0_156_12 (.ZN (n_0_156_11), .A (sps__n74));
INV_X1 i_0_156_11 (.ZN (n_0_156_10), .A (sps__n7));
INV_X1 i_0_156_10 (.ZN (n_0_156_9), .A (sps__n14));
INV_X1 i_0_156_9 (.ZN (n_0_156_8), .A (sps__n85));
INV_X1 i_0_156_8 (.ZN (n_0_156_7), .A (sps__n36));
INV_X1 i_0_156_7 (.ZN (n_0_156_6), .A (address[7]));
INV_X1 i_0_156_6 (.ZN (n_0_156_5), .A (sps__n69));
INV_X1 i_0_156_5 (.ZN (n_0_156_4), .A (sps__n26));
INV_X1 i_0_156_4 (.ZN (n_0_156_3), .A (sps__n42));
INV_X1 i_0_156_3 (.ZN (n_0_156_2), .A (sps__n50));
INV_X1 i_0_156_2 (.ZN (n_0_156_1), .A (sps__n56));
NAND4_X1 i_0_156_1 (.ZN (n_0_156_0), .A1 (n_0_156_26), .A2 (n_0_156_25), .A3 (n_0_156_24), .A4 (data[12]));
NAND2_X1 i_0_156_0 (.ZN (n_0_61), .A1 (n_0_156_19), .A2 (n_0_156_0));
NAND3_X1 i_0_139_36 (.ZN (n_0_60), .A1 (n_0_139_33), .A2 (n_0_139_34), .A3 (n_0_139_35));
NAND2_X1 i_0_139_35 (.ZN (n_0_139_35), .A1 (n_0_139_24), .A2 (\mem[4][12] ));
NAND2_X1 i_0_139_34 (.ZN (n_0_139_34), .A1 (n_0_139_23), .A2 (\mem[4][12] ));
NAND3_X1 i_0_139_33 (.ZN (n_0_139_33), .A1 (n_0_139_26), .A2 (n_0_139_32), .A3 (n_0_139_29));
NOR2_X1 i_0_139_32 (.ZN (n_0_139_32), .A1 (n_0_139_0), .A2 (n_0_139_18));
INV_X1 i_0_139_31 (.ZN (n_0_139_31), .A (n_0_139_18));
INV_X1 i_0_139_30 (.ZN (n_0_139_30), .A (n_0_139_0));
NOR2_X1 i_0_139_29 (.ZN (n_0_139_29), .A1 (n_0_139_5), .A2 (n_0_139_14));
INV_X1 i_0_139_28 (.ZN (n_0_139_28), .A (n_0_139_14));
INV_X1 i_0_139_27 (.ZN (n_0_139_27), .A (n_0_139_5));
INV_X1 i_0_139_26 (.ZN (n_0_139_26), .A (n_0_139_25));
NAND2_X1 i_0_139_25 (.ZN (n_0_139_25), .A1 (n_0_139_10), .A2 (data[12]));
NAND2_X1 i_0_139_24 (.ZN (n_0_139_24), .A1 (n_0_139_30), .A2 (n_0_139_27));
NAND3_X1 i_0_139_23 (.ZN (n_0_139_23), .A1 (n_0_139_31), .A2 (n_0_139_28), .A3 (n_0_139_10));
INV_X1 i_0_139_22 (.ZN (n_0_139_22), .A (sps__n36));
INV_X1 i_0_139_21 (.ZN (n_0_139_21), .A (sps__n9));
INV_X1 i_0_139_20 (.ZN (n_0_139_20), .A (sps__n15));
INV_X1 i_0_139_19 (.ZN (n_0_139_19), .A (sps__n51));
NAND4_X1 i_0_139_18 (.ZN (n_0_139_18), .A1 (n_0_139_22), .A2 (n_0_139_21), .A3 (n_0_139_20), .A4 (n_0_139_19));
INV_X1 i_0_139_17 (.ZN (n_0_139_17), .A (sps__n62));
INV_X1 i_0_139_12 (.ZN (n_0_139_16), .A (sps__n74));
INV_X1 i_0_139_11 (.ZN (n_0_139_15), .A (sps__n86));
NAND4_X1 i_0_139_6 (.ZN (n_0_139_14), .A1 (n_0_139_17), .A2 (n_0_139_16), .A3 (n_0_139_15), .A4 (sps__n2));
INV_X1 i_0_139_5 (.ZN (n_0_139_13), .A (sps__n114));
INV_X1 i_0_139_4 (.ZN (n_0_139_12), .A (sps__n98));
NAND3_X1 i_0_139_1 (.ZN (n_0_139_11), .A1 (n_0_139_13), .A2 (n_0_139_12), .A3 (sps__n123));
INV_X1 i_0_139_0 (.ZN (n_0_139_10), .A (n_0_139_11));
INV_X1 i_0_139_16 (.ZN (n_0_139_9), .A (sps__n68));
INV_X1 i_0_139_15 (.ZN (n_0_139_8), .A (sps__n20));
INV_X1 i_0_139_14 (.ZN (n_0_139_7), .A (sps__n80));
INV_X1 i_0_139_13 (.ZN (n_0_139_6), .A (sps__n103));
NAND4_X1 i_0_139_3 (.ZN (n_0_139_5), .A1 (n_0_139_9), .A2 (n_0_139_8), .A3 (n_0_139_7), .A4 (n_0_139_6));
INV_X1 i_0_139_10 (.ZN (n_0_139_4), .A (sps__n55));
INV_X1 i_0_139_9 (.ZN (n_0_139_3), .A (sps__n28));
INV_X1 i_0_139_8 (.ZN (n_0_139_2), .A (sps__n42));
INV_X1 i_0_139_7 (.ZN (n_0_139_1), .A (sps__n91));
NAND4_X1 i_0_139_2 (.ZN (n_0_139_0), .A1 (n_0_139_4), .A2 (n_0_139_3), .A3 (n_0_139_2), .A4 (n_0_139_1));
NAND3_X1 i_0_122_31 (.ZN (n_0_122_30), .A1 (n_0_122_27), .A2 (n_0_122_28), .A3 (n_0_122_29));
NOR2_X1 i_0_122_30 (.ZN (n_0_122_29), .A1 (n_0_122_13), .A2 (n_0_122_23));
NOR2_X1 i_0_122_29 (.ZN (n_0_122_28), .A1 (n_0_122_22), .A2 (n_0_122_21));
NOR2_X1 i_0_122_28 (.ZN (n_0_122_27), .A1 (n_0_122_17), .A2 (n_0_122_20));
NOR2_X1 i_0_122_27 (.ZN (n_0_122_26), .A1 (n_0_122_17), .A2 (n_0_122_13));
NOR2_X1 i_0_122_26 (.ZN (n_0_122_25), .A1 (n_0_122_20), .A2 (n_0_122_21));
NOR2_X1 i_0_122_25 (.ZN (n_0_122_24), .A1 (n_0_122_22), .A2 (n_0_122_23));
NAND3_X1 i_0_122_24 (.ZN (n_0_122_23), .A1 (n_0_122_4), .A2 (n_0_122_2), .A3 (n_0_122_6));
NAND3_X1 i_0_122_23 (.ZN (n_0_122_22), .A1 (n_0_122_1), .A2 (n_0_122_3), .A3 (n_0_122_5));
NAND3_X1 i_0_122_22 (.ZN (n_0_122_21), .A1 (n_0_122_10), .A2 (n_0_122_8), .A3 (n_0_122_12));
NAND3_X1 i_0_122_21 (.ZN (n_0_122_20), .A1 (n_0_122_7), .A2 (n_0_122_9), .A3 (n_0_122_11));
NAND2_X1 i_0_122_20 (.ZN (n_0_122_19), .A1 (n_0_122_30), .A2 (\mem[5][12] ));
INV_X1 i_0_122_19 (.ZN (n_0_122_18), .A (sps__n114));
NAND4_X1 i_0_122_18 (.ZN (n_0_122_17), .A1 (n_0_122_18), .A2 (sps__n2), .A3 (sps__n123), .A4 (sps__n98));
INV_X1 i_0_122_17 (.ZN (n_0_122_16), .A (sps__n20));
INV_X1 i_0_122_16 (.ZN (n_0_122_15), .A (address[4]));
INV_X1 i_0_122_15 (.ZN (n_0_122_14), .A (sps__n103));
NAND3_X1 i_0_122_14 (.ZN (n_0_122_13), .A1 (n_0_122_16), .A2 (n_0_122_15), .A3 (n_0_122_14));
INV_X1 i_0_122_13 (.ZN (n_0_122_12), .A (RST));
INV_X1 i_0_122_12 (.ZN (n_0_122_11), .A (sps__n74));
INV_X1 i_0_122_11 (.ZN (n_0_122_10), .A (sps__n7));
INV_X1 i_0_122_10 (.ZN (n_0_122_9), .A (sps__n14));
INV_X1 i_0_122_9 (.ZN (n_0_122_8), .A (sps__n85));
INV_X1 i_0_122_8 (.ZN (n_0_122_7), .A (sps__n36));
INV_X1 i_0_122_7 (.ZN (n_0_122_6), .A (sps__n92));
INV_X1 i_0_122_6 (.ZN (n_0_122_5), .A (sps__n69));
INV_X1 i_0_122_5 (.ZN (n_0_122_4), .A (sps__n26));
INV_X1 i_0_122_4 (.ZN (n_0_122_3), .A (sps__n42));
INV_X1 i_0_122_3 (.ZN (n_0_122_2), .A (sps__n50));
INV_X1 i_0_122_2 (.ZN (n_0_122_1), .A (sps__n55));
NAND4_X1 i_0_122_1 (.ZN (n_0_122_0), .A1 (n_0_122_26), .A2 (n_0_122_25), .A3 (n_0_122_24), .A4 (data[12]));
NAND2_X1 i_0_122_0 (.ZN (n_0_59), .A1 (n_0_122_19), .A2 (n_0_122_0));
NAND3_X1 i_0_105_31 (.ZN (n_0_105_30), .A1 (n_0_105_27), .A2 (n_0_105_28), .A3 (n_0_105_29));
NOR2_X1 i_0_105_30 (.ZN (n_0_105_29), .A1 (n_0_105_13), .A2 (n_0_105_23));
NOR2_X1 i_0_105_29 (.ZN (n_0_105_28), .A1 (n_0_105_22), .A2 (n_0_105_21));
NOR2_X1 i_0_105_28 (.ZN (n_0_105_27), .A1 (n_0_105_17), .A2 (n_0_105_20));
NOR2_X1 i_0_105_27 (.ZN (n_0_105_26), .A1 (n_0_105_17), .A2 (n_0_105_13));
NOR2_X1 i_0_105_26 (.ZN (n_0_105_25), .A1 (n_0_105_20), .A2 (n_0_105_21));
NOR2_X1 i_0_105_25 (.ZN (n_0_105_24), .A1 (n_0_105_22), .A2 (n_0_105_23));
NAND3_X1 i_0_105_24 (.ZN (n_0_105_23), .A1 (n_0_105_4), .A2 (n_0_105_2), .A3 (n_0_105_6));
NAND3_X1 i_0_105_23 (.ZN (n_0_105_22), .A1 (n_0_105_1), .A2 (n_0_105_3), .A3 (n_0_105_5));
NAND3_X1 i_0_105_22 (.ZN (n_0_105_21), .A1 (n_0_105_10), .A2 (n_0_105_8), .A3 (n_0_105_12));
NAND3_X1 i_0_105_21 (.ZN (n_0_105_20), .A1 (n_0_105_7), .A2 (n_0_105_9), .A3 (n_0_105_11));
NAND2_X1 i_0_105_20 (.ZN (n_0_105_19), .A1 (n_0_105_30), .A2 (\mem[6][12] ));
INV_X1 i_0_105_19 (.ZN (n_0_105_18), .A (sps__n98));
NAND4_X1 i_0_105_18 (.ZN (n_0_105_17), .A1 (n_0_105_18), .A2 (sps__n2), .A3 (sps__n123), .A4 (sps__n114));
INV_X1 i_0_105_17 (.ZN (n_0_105_16), .A (sps__n19));
INV_X1 i_0_105_16 (.ZN (n_0_105_15), .A (sps__n81));
INV_X1 i_0_105_15 (.ZN (n_0_105_14), .A (sps__n104));
NAND3_X1 i_0_105_14 (.ZN (n_0_105_13), .A1 (n_0_105_16), .A2 (n_0_105_15), .A3 (n_0_105_14));
INV_X1 i_0_105_13 (.ZN (n_0_105_12), .A (sps__n62));
INV_X1 i_0_105_12 (.ZN (n_0_105_11), .A (sps__n74));
INV_X1 i_0_105_11 (.ZN (n_0_105_10), .A (sps__n8));
INV_X1 i_0_105_10 (.ZN (n_0_105_9), .A (sps__n15));
INV_X1 i_0_105_9 (.ZN (n_0_105_8), .A (sps__n86));
INV_X1 i_0_105_8 (.ZN (n_0_105_7), .A (sps__n36));
INV_X1 i_0_105_7 (.ZN (n_0_105_6), .A (sps__n91));
INV_X1 i_0_105_6 (.ZN (n_0_105_5), .A (sps__n68));
INV_X1 i_0_105_5 (.ZN (n_0_105_4), .A (sps__n26));
INV_X1 i_0_105_4 (.ZN (n_0_105_3), .A (sps__n44));
INV_X1 i_0_105_3 (.ZN (n_0_105_2), .A (sps__n50));
INV_X1 i_0_105_2 (.ZN (n_0_105_1), .A (sps__n55));
NAND4_X1 i_0_105_1 (.ZN (n_0_105_0), .A1 (n_0_105_26), .A2 (n_0_105_25), .A3 (n_0_105_24), .A4 (data[12]));
NAND2_X1 i_0_105_0 (.ZN (n_0_58), .A1 (n_0_105_19), .A2 (n_0_105_0));
NAND3_X1 i_0_88_27 (.ZN (n_0_88_26), .A1 (n_0_88_23), .A2 (n_0_88_24), .A3 (n_0_88_25));
NOR2_X1 i_0_88_26 (.ZN (n_0_88_25), .A1 (n_0_88_17), .A2 (n_0_88_13));
NOR2_X1 i_0_88_25 (.ZN (n_0_88_24), .A1 (n_0_88_19), .A2 (n_0_88_20));
NOR2_X1 i_0_88_24 (.ZN (n_0_88_23), .A1 (n_0_88_21), .A2 (n_0_88_22));
NAND3_X1 i_0_88_23 (.ZN (n_0_88_22), .A1 (n_0_88_4), .A2 (n_0_88_2), .A3 (n_0_88_6));
NAND3_X1 i_0_88_22 (.ZN (n_0_88_21), .A1 (n_0_88_1), .A2 (n_0_88_3), .A3 (n_0_88_5));
NAND3_X1 i_0_88_21 (.ZN (n_0_88_20), .A1 (n_0_88_10), .A2 (n_0_88_8), .A3 (n_0_88_12));
NAND3_X1 i_0_88_20 (.ZN (n_0_88_19), .A1 (n_0_88_7), .A2 (n_0_88_9), .A3 (n_0_88_11));
NAND2_X1 i_0_88_19 (.ZN (n_0_88_18), .A1 (n_0_88_26), .A2 (\mem[7][12] ));
NAND4_X1 i_0_88_18 (.ZN (n_0_88_17), .A1 (sps__n2), .A2 (sps__n123), .A3 (sps__n114), .A4 (sps__n98));
INV_X1 i_0_88_17 (.ZN (n_0_88_16), .A (sps__n20));
INV_X1 i_0_88_16 (.ZN (n_0_88_15), .A (sps__n80));
INV_X1 i_0_88_15 (.ZN (n_0_88_14), .A (sps__n104));
NAND3_X1 i_0_88_14 (.ZN (n_0_88_13), .A1 (n_0_88_16), .A2 (n_0_88_15), .A3 (n_0_88_14));
INV_X1 i_0_88_13 (.ZN (n_0_88_12), .A (RST));
INV_X1 i_0_88_12 (.ZN (n_0_88_11), .A (sps__n74));
INV_X1 i_0_88_11 (.ZN (n_0_88_10), .A (sps__n7));
INV_X1 i_0_88_10 (.ZN (n_0_88_9), .A (sps__n14));
INV_X1 i_0_88_9 (.ZN (n_0_88_8), .A (sps__n85));
INV_X1 i_0_88_8 (.ZN (n_0_88_7), .A (sps__n36));
INV_X1 i_0_88_7 (.ZN (n_0_88_6), .A (sps__n91));
INV_X1 i_0_88_6 (.ZN (n_0_88_5), .A (sps__n69));
INV_X1 i_0_88_5 (.ZN (n_0_88_4), .A (sps__n26));
INV_X1 i_0_88_4 (.ZN (n_0_88_3), .A (sps__n42));
INV_X1 i_0_88_3 (.ZN (n_0_88_2), .A (sps__n50));
INV_X1 i_0_88_2 (.ZN (n_0_88_1), .A (sps__n56));
NAND4_X1 i_0_88_1 (.ZN (n_0_88_0), .A1 (n_0_88_25), .A2 (n_0_88_24), .A3 (n_0_88_23), .A4 (data[12]));
NAND2_X1 i_0_88_0 (.ZN (n_0_57), .A1 (n_0_88_18), .A2 (n_0_88_0));
NAND3_X1 i_0_71_35 (.ZN (n_0_56), .A1 (n_0_71_32), .A2 (n_0_71_33), .A3 (n_0_71_34));
NAND2_X1 i_0_71_34 (.ZN (n_0_71_34), .A1 (n_0_71_23), .A2 (\mem[8][12] ));
NAND3_X1 i_0_71_29 (.ZN (n_0_71_33), .A1 (n_0_71_26), .A2 (n_0_71_31), .A3 (n_0_71_28));
NAND2_X1 i_0_71_28 (.ZN (n_0_71_32), .A1 (n_0_71_27), .A2 (\mem[8][12] ));
NOR2_X1 i_0_71_24 (.ZN (n_0_71_31), .A1 (n_0_71_18), .A2 (n_0_71_0));
INV_X1 i_0_71_23 (.ZN (n_0_71_30), .A (n_0_71_0));
INV_X1 i_0_71_22 (.ZN (n_0_71_29), .A (n_0_71_18));
INV_X1 i_0_71_21 (.ZN (n_0_71_28), .A (n_0_71_5));
NAND3_X1 i_0_71_20 (.ZN (n_0_71_27), .A1 (n_0_71_28), .A2 (n_0_71_30), .A3 (n_0_71_9));
NOR2_X1 i_0_71_19 (.ZN (n_0_71_26), .A1 (n_0_71_14), .A2 (n_0_71_24));
INV_X1 i_0_71_18 (.ZN (n_0_71_25), .A (n_0_71_14));
NAND2_X1 i_0_71_17 (.ZN (n_0_71_24), .A1 (n_0_71_9), .A2 (data[12]));
NAND2_X1 i_0_71_16 (.ZN (n_0_71_23), .A1 (n_0_71_29), .A2 (n_0_71_25));
INV_X1 i_0_71_33 (.ZN (n_0_71_22), .A (sps__n36));
INV_X1 i_0_71_32 (.ZN (n_0_71_21), .A (sps__n9));
INV_X1 i_0_71_31 (.ZN (n_0_71_20), .A (sps__n14));
INV_X1 i_0_71_30 (.ZN (n_0_71_19), .A (sps__n51));
NAND4_X1 i_0_71_3 (.ZN (n_0_71_18), .A1 (n_0_71_22), .A2 (n_0_71_21), .A3 (n_0_71_20), .A4 (n_0_71_19));
INV_X1 i_0_71_27 (.ZN (n_0_71_17), .A (sps__n62));
INV_X1 i_0_71_26 (.ZN (n_0_71_16), .A (sps__n74));
INV_X1 i_0_71_25 (.ZN (n_0_71_15), .A (sps__n86));
NAND4_X1 i_0_71_8 (.ZN (n_0_71_14), .A1 (n_0_71_17), .A2 (n_0_71_16), .A3 (n_0_71_15), .A4 (sps__n2));
INV_X1 i_0_71_15 (.ZN (n_0_71_13), .A (sps__n123));
INV_X1 i_0_71_14 (.ZN (n_0_71_12), .A (sps__n114));
INV_X1 i_0_71_13 (.ZN (n_0_71_11), .A (sps__n98));
NAND3_X1 i_0_71_12 (.ZN (n_0_71_10), .A1 (n_0_71_13), .A2 (n_0_71_12), .A3 (n_0_71_11));
INV_X1 i_0_71_11 (.ZN (n_0_71_9), .A (n_0_71_10));
INV_X1 i_0_71_10 (.ZN (n_0_71_8), .A (sps__n68));
INV_X1 i_0_71_9 (.ZN (n_0_71_7), .A (sps__n20));
INV_X1 i_0_71_7 (.ZN (n_0_71_6), .A (sps__n80));
NAND4_X1 i_0_71_6 (.ZN (n_0_71_5), .A1 (n_0_71_8), .A2 (n_0_71_7), .A3 (n_0_71_6), .A4 (sps__n103));
INV_X1 i_0_71_5 (.ZN (n_0_71_4), .A (sps__n55));
INV_X1 i_0_71_4 (.ZN (n_0_71_3), .A (address[9]));
INV_X1 i_0_71_2 (.ZN (n_0_71_2), .A (sps__n42));
INV_X1 i_0_71_1 (.ZN (n_0_71_1), .A (sps__n92));
NAND4_X1 i_0_71_0 (.ZN (n_0_71_0), .A1 (n_0_71_4), .A2 (n_0_71_3), .A3 (n_0_71_2), .A4 (n_0_71_1));
NOR2_X1 i_0_54_34 (.ZN (n_0_54_33), .A1 (n_0_54_19), .A2 (n_0_54_0));
INV_X1 i_0_54_33 (.ZN (n_0_54_32), .A (n_0_54_0));
INV_X1 i_0_54_28 (.ZN (n_0_54_31), .A (n_0_54_19));
NAND2_X1 i_0_54_27 (.ZN (n_0_54_30), .A1 (n_0_54_29), .A2 (\mem[9][12] ));
NAND3_X1 i_0_54_23 (.ZN (n_0_54_29), .A1 (n_0_54_5), .A2 (n_0_54_32), .A3 (n_0_54_10));
NAND3_X1 i_0_54_22 (.ZN (n_0_54_28), .A1 (n_0_54_27), .A2 (n_0_54_33), .A3 (n_0_54_14));
NOR2_X1 i_0_54_21 (.ZN (n_0_54_27), .A1 (n_0_54_6), .A2 (n_0_54_26));
NAND2_X1 i_0_54_20 (.ZN (n_0_54_26), .A1 (n_0_54_10), .A2 (data[12]));
NAND2_X1 i_0_54_19 (.ZN (n_0_54_25), .A1 (n_0_54_31), .A2 (n_0_54_14));
NAND3_X1 i_0_54_18 (.ZN (n_0_55), .A1 (n_0_54_28), .A2 (n_0_54_30), .A3 (n_0_54_24));
NAND2_X1 i_0_54_17 (.ZN (n_0_54_24), .A1 (n_0_54_25), .A2 (\mem[9][12] ));
INV_X1 i_0_54_32 (.ZN (n_0_54_23), .A (sps__n36));
INV_X1 i_0_54_31 (.ZN (n_0_54_22), .A (sps__n7));
INV_X1 i_0_54_30 (.ZN (n_0_54_21), .A (sps__n14));
INV_X1 i_0_54_29 (.ZN (n_0_54_20), .A (sps__n50));
NAND4_X1 i_0_54_3 (.ZN (n_0_54_19), .A1 (n_0_54_23), .A2 (n_0_54_22), .A3 (n_0_54_21), .A4 (n_0_54_20));
INV_X1 i_0_54_26 (.ZN (n_0_54_18), .A (RST));
INV_X1 i_0_54_25 (.ZN (n_0_54_17), .A (sps__n74));
INV_X1 i_0_54_24 (.ZN (n_0_54_16), .A (sps__n85));
NAND4_X1 i_0_54_6 (.ZN (n_0_54_15), .A1 (n_0_54_18), .A2 (n_0_54_17), .A3 (n_0_54_16), .A4 (sps__n2));
INV_X1 i_0_54_16 (.ZN (n_0_54_14), .A (n_0_54_15));
INV_X1 i_0_54_15 (.ZN (n_0_54_13), .A (sps__n123));
INV_X1 i_0_54_14 (.ZN (n_0_54_12), .A (sps__n114));
NAND3_X1 i_0_54_13 (.ZN (n_0_54_11), .A1 (n_0_54_13), .A2 (n_0_54_12), .A3 (sps__n98));
INV_X1 i_0_54_12 (.ZN (n_0_54_10), .A (n_0_54_11));
INV_X1 i_0_54_11 (.ZN (n_0_54_9), .A (sps__n69));
INV_X1 i_0_54_10 (.ZN (n_0_54_8), .A (sps__n20));
INV_X1 i_0_54_9 (.ZN (n_0_54_7), .A (address[4]));
NAND4_X1 i_0_54_8 (.ZN (n_0_54_6), .A1 (n_0_54_9), .A2 (n_0_54_8), .A3 (n_0_54_7), .A4 (sps__n103));
INV_X1 i_0_54_7 (.ZN (n_0_54_5), .A (n_0_54_6));
INV_X1 i_0_54_5 (.ZN (n_0_54_4), .A (sps__n56));
INV_X1 i_0_54_4 (.ZN (n_0_54_3), .A (sps__n26));
INV_X1 i_0_54_2 (.ZN (n_0_54_2), .A (sps__n42));
INV_X1 i_0_54_1 (.ZN (n_0_54_1), .A (address[7]));
NAND4_X1 i_0_54_0 (.ZN (n_0_54_0), .A1 (n_0_54_4), .A2 (n_0_54_3), .A3 (n_0_54_2), .A4 (n_0_54_1));
NOR2_X1 i_0_37_34 (.ZN (n_0_37_33), .A1 (n_0_37_19), .A2 (n_0_37_0));
INV_X1 i_0_37_33 (.ZN (n_0_37_32), .A (n_0_37_0));
INV_X1 i_0_37_28 (.ZN (n_0_37_31), .A (n_0_37_19));
NAND2_X1 i_0_37_27 (.ZN (n_0_37_30), .A1 (n_0_37_29), .A2 (\mem[10][12] ));
NAND3_X1 i_0_37_23 (.ZN (n_0_37_29), .A1 (n_0_37_5), .A2 (n_0_37_32), .A3 (n_0_37_10));
NAND3_X1 i_0_37_22 (.ZN (n_0_37_28), .A1 (n_0_37_27), .A2 (n_0_37_33), .A3 (n_0_37_14));
NOR2_X1 i_0_37_21 (.ZN (n_0_37_27), .A1 (n_0_37_6), .A2 (n_0_37_26));
NAND2_X1 i_0_37_20 (.ZN (n_0_37_26), .A1 (n_0_37_10), .A2 (data[12]));
NAND2_X1 i_0_37_19 (.ZN (n_0_37_25), .A1 (n_0_37_31), .A2 (n_0_37_14));
NAND3_X1 i_0_37_18 (.ZN (n_0_54), .A1 (n_0_37_28), .A2 (n_0_37_30), .A3 (n_0_37_24));
NAND2_X1 i_0_37_17 (.ZN (n_0_37_24), .A1 (n_0_37_25), .A2 (\mem[10][12] ));
INV_X1 i_0_37_32 (.ZN (n_0_37_23), .A (sps__n36));
INV_X1 i_0_37_31 (.ZN (n_0_37_22), .A (sps__n7));
INV_X1 i_0_37_30 (.ZN (n_0_37_21), .A (sps__n14));
INV_X1 i_0_37_29 (.ZN (n_0_37_20), .A (sps__n50));
NAND4_X1 i_0_37_3 (.ZN (n_0_37_19), .A1 (n_0_37_23), .A2 (n_0_37_22), .A3 (n_0_37_21), .A4 (n_0_37_20));
INV_X1 i_0_37_26 (.ZN (n_0_37_18), .A (sps__n61));
INV_X1 i_0_37_25 (.ZN (n_0_37_17), .A (sps__n74));
INV_X1 i_0_37_24 (.ZN (n_0_37_16), .A (sps__n85));
NAND4_X1 i_0_37_6 (.ZN (n_0_37_15), .A1 (n_0_37_18), .A2 (n_0_37_17), .A3 (n_0_37_16), .A4 (sps__n2));
INV_X1 i_0_37_16 (.ZN (n_0_37_14), .A (n_0_37_15));
INV_X1 i_0_37_15 (.ZN (n_0_37_13), .A (sps__n121));
INV_X1 i_0_37_14 (.ZN (n_0_37_12), .A (sps__n97));
NAND3_X1 i_0_37_13 (.ZN (n_0_37_11), .A1 (n_0_37_13), .A2 (n_0_37_12), .A3 (sps__n114));
INV_X1 i_0_37_12 (.ZN (n_0_37_10), .A (n_0_37_11));
INV_X1 i_0_37_11 (.ZN (n_0_37_9), .A (sps__n68));
INV_X1 i_0_37_10 (.ZN (n_0_37_8), .A (sps__n20));
INV_X1 i_0_37_9 (.ZN (n_0_37_7), .A (sps__n80));
NAND4_X1 i_0_37_8 (.ZN (n_0_37_6), .A1 (n_0_37_9), .A2 (n_0_37_8), .A3 (n_0_37_7), .A4 (sps__n104));
INV_X1 i_0_37_7 (.ZN (n_0_37_5), .A (n_0_37_6));
INV_X1 i_0_37_5 (.ZN (n_0_37_4), .A (sps__n55));
INV_X1 i_0_37_4 (.ZN (n_0_37_3), .A (sps__n26));
INV_X1 i_0_37_2 (.ZN (n_0_37_2), .A (sps__n44));
INV_X1 i_0_37_1 (.ZN (n_0_37_1), .A (sps__n91));
NAND4_X1 i_0_37_0 (.ZN (n_0_37_0), .A1 (n_0_37_4), .A2 (n_0_37_3), .A3 (n_0_37_2), .A4 (n_0_37_1));
NAND3_X1 i_0_20_37 (.ZN (n_0_53), .A1 (n_0_20_34), .A2 (n_0_20_35), .A3 (n_0_20_36));
NAND2_X1 i_0_20_36 (.ZN (n_0_20_36), .A1 (n_0_20_25), .A2 (\mem[0][13] ));
NAND3_X1 i_0_20_35 (.ZN (n_0_20_35), .A1 (n_0_20_27), .A2 (n_0_20_33), .A3 (n_0_20_30));
NAND2_X1 i_0_20_34 (.ZN (n_0_20_34), .A1 (n_0_20_24), .A2 (\mem[0][13] ));
NOR2_X1 i_0_20_33 (.ZN (n_0_20_33), .A1 (n_0_20_0), .A2 (n_0_20_19));
INV_X1 i_0_20_32 (.ZN (n_0_20_32), .A (n_0_20_19));
INV_X1 i_0_20_31 (.ZN (n_0_20_31), .A (n_0_20_0));
NOR2_X1 i_0_20_30 (.ZN (n_0_20_30), .A1 (n_0_20_5), .A2 (n_0_20_15));
INV_X1 i_0_20_29 (.ZN (n_0_20_29), .A (n_0_20_15));
INV_X1 i_0_20_28 (.ZN (n_0_20_28), .A (n_0_20_5));
INV_X1 i_0_20_27 (.ZN (n_0_20_27), .A (n_0_20_26));
NAND2_X1 i_0_20_26 (.ZN (n_0_20_26), .A1 (n_0_20_10), .A2 (data[13]));
NAND2_X1 i_0_20_25 (.ZN (n_0_20_25), .A1 (n_0_20_31), .A2 (n_0_20_28));
NAND3_X1 i_0_20_24 (.ZN (n_0_20_24), .A1 (n_0_20_32), .A2 (n_0_20_29), .A3 (n_0_20_10));
INV_X1 i_0_20_23 (.ZN (n_0_20_23), .A (sps__n34));
INV_X1 i_0_20_22 (.ZN (n_0_20_22), .A (sps__n9));
INV_X1 i_0_20_21 (.ZN (n_0_20_21), .A (sps__n15));
INV_X1 i_0_20_20 (.ZN (n_0_20_20), .A (sps__n51));
NAND4_X1 i_0_20_19 (.ZN (n_0_20_19), .A1 (n_0_20_23), .A2 (n_0_20_22), .A3 (n_0_20_21), .A4 (n_0_20_20));
INV_X1 i_0_20_18 (.ZN (n_0_20_18), .A (sps__n62));
INV_X1 i_0_20_17 (.ZN (n_0_20_17), .A (sps__n74));
INV_X1 i_0_20_12 (.ZN (n_0_20_16), .A (sps__n86));
NAND4_X1 i_0_20_11 (.ZN (n_0_20_15), .A1 (n_0_20_18), .A2 (n_0_20_17), .A3 (n_0_20_16), .A4 (sps__n3));
INV_X1 i_0_20_6 (.ZN (n_0_20_14), .A (sps__n122));
INV_X1 i_0_20_5 (.ZN (n_0_20_13), .A (sps__n112));
INV_X1 i_0_20_4 (.ZN (n_0_20_12), .A (sps__n99));
NAND3_X1 i_0_20_1 (.ZN (n_0_20_11), .A1 (n_0_20_14), .A2 (n_0_20_13), .A3 (n_0_20_12));
INV_X1 i_0_20_0 (.ZN (n_0_20_10), .A (n_0_20_11));
INV_X1 i_0_20_16 (.ZN (n_0_20_9), .A (sps__n68));
INV_X1 i_0_20_15 (.ZN (n_0_20_8), .A (sps__n19));
INV_X1 i_0_20_14 (.ZN (n_0_20_7), .A (sps__n81));
INV_X1 i_0_20_13 (.ZN (n_0_20_6), .A (sps__n104));
NAND4_X1 i_0_20_3 (.ZN (n_0_20_5), .A1 (n_0_20_9), .A2 (n_0_20_8), .A3 (n_0_20_7), .A4 (n_0_20_6));
INV_X1 i_0_20_10 (.ZN (n_0_20_4), .A (sps__n55));
INV_X1 i_0_20_9 (.ZN (n_0_20_3), .A (sps__n28));
INV_X1 i_0_20_8 (.ZN (n_0_20_2), .A (sps__n43));
INV_X1 i_0_20_7 (.ZN (n_0_20_1), .A (sps__n92));
NAND4_X1 i_0_20_2 (.ZN (n_0_20_0), .A1 (n_0_20_4), .A2 (n_0_20_3), .A3 (n_0_20_2), .A4 (n_0_20_1));
NAND3_X1 i_0_50_36 (.ZN (n_0_52), .A1 (n_0_50_33), .A2 (n_0_50_34), .A3 (n_0_50_35));
NAND2_X1 i_0_50_35 (.ZN (n_0_50_35), .A1 (n_0_50_24), .A2 (\mem[1][13] ));
NAND2_X1 i_0_50_34 (.ZN (n_0_50_34), .A1 (n_0_50_23), .A2 (\mem[1][13] ));
NAND3_X1 i_0_50_33 (.ZN (n_0_50_33), .A1 (n_0_50_26), .A2 (n_0_50_32), .A3 (n_0_50_29));
NOR2_X1 i_0_50_32 (.ZN (n_0_50_32), .A1 (n_0_50_0), .A2 (n_0_50_18));
INV_X1 i_0_50_31 (.ZN (n_0_50_31), .A (n_0_50_18));
INV_X1 i_0_50_30 (.ZN (n_0_50_30), .A (n_0_50_0));
NOR2_X1 i_0_50_29 (.ZN (n_0_50_29), .A1 (n_0_50_5), .A2 (n_0_50_14));
INV_X1 i_0_50_28 (.ZN (n_0_50_28), .A (n_0_50_14));
INV_X1 i_0_50_27 (.ZN (n_0_50_27), .A (n_0_50_5));
INV_X1 i_0_50_26 (.ZN (n_0_50_26), .A (n_0_50_25));
NAND2_X1 i_0_50_25 (.ZN (n_0_50_25), .A1 (n_0_50_10), .A2 (data[13]));
NAND2_X1 i_0_50_24 (.ZN (n_0_50_24), .A1 (n_0_50_30), .A2 (n_0_50_27));
NAND3_X1 i_0_50_23 (.ZN (n_0_50_23), .A1 (n_0_50_31), .A2 (n_0_50_28), .A3 (n_0_50_10));
INV_X1 i_0_50_22 (.ZN (n_0_50_22), .A (sps__n35));
INV_X1 i_0_50_21 (.ZN (n_0_50_21), .A (sps__n8));
INV_X1 i_0_50_20 (.ZN (n_0_50_20), .A (sps__n13));
INV_X1 i_0_50_19 (.ZN (n_0_50_19), .A (sps__n49));
NAND4_X1 i_0_50_18 (.ZN (n_0_50_18), .A1 (n_0_50_22), .A2 (n_0_50_21), .A3 (n_0_50_20), .A4 (n_0_50_19));
INV_X1 i_0_50_17 (.ZN (n_0_50_17), .A (sps__n63));
INV_X1 i_0_50_12 (.ZN (n_0_50_16), .A (sps__n74));
INV_X1 i_0_50_11 (.ZN (n_0_50_15), .A (sps__n87));
NAND4_X1 i_0_50_6 (.ZN (n_0_50_14), .A1 (n_0_50_17), .A2 (n_0_50_16), .A3 (n_0_50_15), .A4 (sps__n1));
INV_X1 i_0_50_5 (.ZN (n_0_50_13), .A (sps__n121));
INV_X1 i_0_50_4 (.ZN (n_0_50_12), .A (sps__n112));
NAND3_X1 i_0_50_1 (.ZN (n_0_50_11), .A1 (n_0_50_13), .A2 (n_0_50_12), .A3 (sps__n97));
INV_X1 i_0_50_0 (.ZN (n_0_50_10), .A (n_0_50_11));
INV_X1 i_0_50_16 (.ZN (n_0_50_9), .A (sps__n68));
INV_X1 i_0_50_15 (.ZN (n_0_50_8), .A (sps__n21));
INV_X1 i_0_50_14 (.ZN (n_0_50_7), .A (sps__n80));
INV_X1 i_0_50_13 (.ZN (n_0_50_6), .A (sps__n103));
NAND4_X1 i_0_50_3 (.ZN (n_0_50_5), .A1 (n_0_50_9), .A2 (n_0_50_8), .A3 (n_0_50_7), .A4 (n_0_50_6));
INV_X1 i_0_50_10 (.ZN (n_0_50_4), .A (sps__n57));
INV_X1 i_0_50_9 (.ZN (n_0_50_3), .A (sps__n26));
INV_X1 i_0_50_8 (.ZN (n_0_50_2), .A (sps__n44));
INV_X1 i_0_50_7 (.ZN (n_0_50_1), .A (sps__n91));
NAND4_X1 i_0_50_2 (.ZN (n_0_50_0), .A1 (n_0_50_4), .A2 (n_0_50_3), .A3 (n_0_50_2), .A4 (n_0_50_1));
NAND3_X1 i_0_172_36 (.ZN (n_0_51), .A1 (n_0_172_33), .A2 (n_0_172_34), .A3 (n_0_172_35));
NAND2_X1 i_0_172_35 (.ZN (n_0_172_35), .A1 (n_0_172_24), .A2 (\mem[2][13] ));
NAND2_X1 i_0_172_34 (.ZN (n_0_172_34), .A1 (n_0_172_23), .A2 (\mem[2][13] ));
NAND3_X1 i_0_172_33 (.ZN (n_0_172_33), .A1 (n_0_172_26), .A2 (n_0_172_32), .A3 (n_0_172_29));
NOR2_X1 i_0_172_32 (.ZN (n_0_172_32), .A1 (n_0_172_0), .A2 (n_0_172_18));
INV_X1 i_0_172_31 (.ZN (n_0_172_31), .A (n_0_172_18));
INV_X1 i_0_172_30 (.ZN (n_0_172_30), .A (n_0_172_0));
NOR2_X1 i_0_172_29 (.ZN (n_0_172_29), .A1 (n_0_172_5), .A2 (n_0_172_14));
INV_X1 i_0_172_28 (.ZN (n_0_172_28), .A (n_0_172_14));
INV_X1 i_0_172_27 (.ZN (n_0_172_27), .A (n_0_172_5));
INV_X1 i_0_172_26 (.ZN (n_0_172_26), .A (n_0_172_25));
NAND2_X1 i_0_172_25 (.ZN (n_0_172_25), .A1 (n_0_172_10), .A2 (data[13]));
NAND2_X1 i_0_172_24 (.ZN (n_0_172_24), .A1 (n_0_172_30), .A2 (n_0_172_27));
NAND3_X1 i_0_172_23 (.ZN (n_0_172_23), .A1 (n_0_172_31), .A2 (n_0_172_28), .A3 (n_0_172_10));
INV_X1 i_0_172_22 (.ZN (n_0_172_22), .A (sps__n36));
INV_X1 i_0_172_21 (.ZN (n_0_172_21), .A (sps__n8));
INV_X1 i_0_172_20 (.ZN (n_0_172_20), .A (sps__n15));
INV_X1 i_0_172_19 (.ZN (n_0_172_19), .A (sps__n50));
NAND4_X1 i_0_172_18 (.ZN (n_0_172_18), .A1 (n_0_172_22), .A2 (n_0_172_21), .A3 (n_0_172_20), .A4 (n_0_172_19));
INV_X1 i_0_172_17 (.ZN (n_0_172_17), .A (sps__n62));
INV_X1 i_0_172_12 (.ZN (n_0_172_16), .A (sps__n74));
INV_X1 i_0_172_11 (.ZN (n_0_172_15), .A (sps__n86));
NAND4_X1 i_0_172_6 (.ZN (n_0_172_14), .A1 (n_0_172_17), .A2 (n_0_172_16), .A3 (n_0_172_15), .A4 (sps__n2));
INV_X1 i_0_172_5 (.ZN (n_0_172_13), .A (sps__n121));
INV_X1 i_0_172_4 (.ZN (n_0_172_12), .A (sps__n99));
NAND3_X1 i_0_172_1 (.ZN (n_0_172_11), .A1 (n_0_172_13), .A2 (n_0_172_12), .A3 (sps__n112));
INV_X1 i_0_172_0 (.ZN (n_0_172_10), .A (n_0_172_11));
INV_X1 i_0_172_16 (.ZN (n_0_172_9), .A (sps__n68));
INV_X1 i_0_172_15 (.ZN (n_0_172_8), .A (sps__n19));
INV_X1 i_0_172_14 (.ZN (n_0_172_7), .A (sps__n81));
INV_X1 i_0_172_13 (.ZN (n_0_172_6), .A (sps__n104));
NAND4_X1 i_0_172_3 (.ZN (n_0_172_5), .A1 (n_0_172_9), .A2 (n_0_172_8), .A3 (n_0_172_7), .A4 (n_0_172_6));
INV_X1 i_0_172_10 (.ZN (n_0_172_4), .A (sps__n55));
INV_X1 i_0_172_9 (.ZN (n_0_172_3), .A (sps__n28));
INV_X1 i_0_172_8 (.ZN (n_0_172_2), .A (sps__n42));
INV_X1 i_0_172_7 (.ZN (n_0_172_1), .A (sps__n91));
NAND4_X1 i_0_172_2 (.ZN (n_0_172_0), .A1 (n_0_172_4), .A2 (n_0_172_3), .A3 (n_0_172_2), .A4 (n_0_172_1));
NAND3_X1 i_0_155_31 (.ZN (n_0_155_30), .A1 (n_0_155_27), .A2 (n_0_155_28), .A3 (n_0_155_29));
NOR2_X1 i_0_155_30 (.ZN (n_0_155_29), .A1 (n_0_155_13), .A2 (n_0_155_23));
NOR2_X1 i_0_155_29 (.ZN (n_0_155_28), .A1 (n_0_155_22), .A2 (n_0_155_21));
NOR2_X1 i_0_155_28 (.ZN (n_0_155_27), .A1 (n_0_155_17), .A2 (n_0_155_20));
NOR2_X1 i_0_155_27 (.ZN (n_0_155_26), .A1 (n_0_155_17), .A2 (n_0_155_13));
NOR2_X1 i_0_155_26 (.ZN (n_0_155_25), .A1 (n_0_155_20), .A2 (n_0_155_21));
NOR2_X1 i_0_155_25 (.ZN (n_0_155_24), .A1 (n_0_155_22), .A2 (n_0_155_23));
NAND3_X1 i_0_155_24 (.ZN (n_0_155_23), .A1 (n_0_155_4), .A2 (n_0_155_2), .A3 (n_0_155_6));
NAND3_X1 i_0_155_23 (.ZN (n_0_155_22), .A1 (n_0_155_1), .A2 (n_0_155_3), .A3 (n_0_155_5));
NAND3_X1 i_0_155_22 (.ZN (n_0_155_21), .A1 (n_0_155_10), .A2 (n_0_155_8), .A3 (n_0_155_12));
NAND3_X1 i_0_155_21 (.ZN (n_0_155_20), .A1 (n_0_155_7), .A2 (n_0_155_9), .A3 (n_0_155_11));
NAND2_X1 i_0_155_20 (.ZN (n_0_155_19), .A1 (n_0_155_30), .A2 (\mem[3][13] ));
INV_X1 i_0_155_19 (.ZN (n_0_155_18), .A (sps__n121));
NAND4_X1 i_0_155_18 (.ZN (n_0_155_17), .A1 (n_0_155_18), .A2 (sps__n1), .A3 (sps__n113), .A4 (sps__n97));
INV_X1 i_0_155_17 (.ZN (n_0_155_16), .A (sps__n21));
INV_X1 i_0_155_16 (.ZN (n_0_155_15), .A (sps__n80));
INV_X1 i_0_155_15 (.ZN (n_0_155_14), .A (sps__n103));
NAND3_X1 i_0_155_14 (.ZN (n_0_155_13), .A1 (n_0_155_16), .A2 (n_0_155_15), .A3 (n_0_155_14));
INV_X1 i_0_155_13 (.ZN (n_0_155_12), .A (sps__n61));
INV_X1 i_0_155_12 (.ZN (n_0_155_11), .A (sps__n74));
INV_X1 i_0_155_11 (.ZN (n_0_155_10), .A (sps__n7));
INV_X1 i_0_155_10 (.ZN (n_0_155_9), .A (sps__n13));
INV_X1 i_0_155_9 (.ZN (n_0_155_8), .A (sps__n87));
INV_X1 i_0_155_8 (.ZN (n_0_155_7), .A (sps__n36));
INV_X1 i_0_155_7 (.ZN (n_0_155_6), .A (sps__n91));
INV_X1 i_0_155_6 (.ZN (n_0_155_5), .A (sps__n69));
INV_X1 i_0_155_5 (.ZN (n_0_155_4), .A (sps__n27));
INV_X1 i_0_155_4 (.ZN (n_0_155_3), .A (sps__n41));
INV_X1 i_0_155_3 (.ZN (n_0_155_2), .A (sps__n49));
INV_X1 i_0_155_2 (.ZN (n_0_155_1), .A (sps__n56));
NAND4_X1 i_0_155_1 (.ZN (n_0_155_0), .A1 (n_0_155_26), .A2 (n_0_155_25), .A3 (n_0_155_24), .A4 (data[13]));
NAND2_X1 i_0_155_0 (.ZN (n_0_50), .A1 (n_0_155_19), .A2 (n_0_155_0));
NAND3_X1 i_0_138_36 (.ZN (n_0_47), .A1 (n_0_138_33), .A2 (n_0_138_34), .A3 (n_0_138_35));
NAND2_X1 i_0_138_35 (.ZN (n_0_138_35), .A1 (n_0_138_24), .A2 (\mem[4][13] ));
NAND2_X1 i_0_138_34 (.ZN (n_0_138_34), .A1 (n_0_138_23), .A2 (\mem[4][13] ));
NAND3_X1 i_0_138_33 (.ZN (n_0_138_33), .A1 (n_0_138_26), .A2 (n_0_138_32), .A3 (n_0_138_29));
NOR2_X1 i_0_138_32 (.ZN (n_0_138_32), .A1 (n_0_138_0), .A2 (n_0_138_18));
INV_X1 i_0_138_31 (.ZN (n_0_138_31), .A (n_0_138_18));
INV_X1 i_0_138_30 (.ZN (n_0_138_30), .A (n_0_138_0));
NOR2_X1 i_0_138_29 (.ZN (n_0_138_29), .A1 (n_0_138_5), .A2 (n_0_138_14));
INV_X1 i_0_138_28 (.ZN (n_0_138_28), .A (n_0_138_14));
INV_X1 i_0_138_27 (.ZN (n_0_138_27), .A (n_0_138_5));
INV_X1 i_0_138_26 (.ZN (n_0_138_26), .A (n_0_138_25));
NAND2_X1 i_0_138_25 (.ZN (n_0_138_25), .A1 (n_0_138_10), .A2 (data[13]));
NAND2_X1 i_0_138_24 (.ZN (n_0_138_24), .A1 (n_0_138_30), .A2 (n_0_138_27));
NAND3_X1 i_0_138_23 (.ZN (n_0_138_23), .A1 (n_0_138_31), .A2 (n_0_138_28), .A3 (n_0_138_10));
INV_X1 i_0_138_22 (.ZN (n_0_138_22), .A (address[14]));
INV_X1 i_0_138_21 (.ZN (n_0_138_21), .A (sps__n9));
INV_X1 i_0_138_20 (.ZN (n_0_138_20), .A (sps__n15));
INV_X1 i_0_138_19 (.ZN (n_0_138_19), .A (sps__n51));
NAND4_X1 i_0_138_18 (.ZN (n_0_138_18), .A1 (n_0_138_22), .A2 (n_0_138_21), .A3 (n_0_138_20), .A4 (n_0_138_19));
INV_X1 i_0_138_17 (.ZN (n_0_138_17), .A (sps__n62));
INV_X1 i_0_138_12 (.ZN (n_0_138_16), .A (sps__n75));
INV_X1 i_0_138_11 (.ZN (n_0_138_15), .A (sps__n86));
NAND4_X1 i_0_138_6 (.ZN (n_0_138_14), .A1 (n_0_138_17), .A2 (n_0_138_16), .A3 (n_0_138_15), .A4 (sps__n2));
INV_X1 i_0_138_5 (.ZN (n_0_138_13), .A (sps__n112));
INV_X1 i_0_138_4 (.ZN (n_0_138_12), .A (sps__n99));
NAND3_X1 i_0_138_1 (.ZN (n_0_138_11), .A1 (n_0_138_13), .A2 (n_0_138_12), .A3 (sps__n121));
INV_X1 i_0_138_0 (.ZN (n_0_138_10), .A (n_0_138_11));
INV_X1 i_0_138_16 (.ZN (n_0_138_9), .A (sps__n68));
INV_X1 i_0_138_15 (.ZN (n_0_138_8), .A (sps__n19));
INV_X1 i_0_138_14 (.ZN (n_0_138_7), .A (sps__n81));
INV_X1 i_0_138_13 (.ZN (n_0_138_6), .A (sps__n105));
NAND4_X1 i_0_138_3 (.ZN (n_0_138_5), .A1 (n_0_138_9), .A2 (n_0_138_8), .A3 (n_0_138_7), .A4 (n_0_138_6));
INV_X1 i_0_138_10 (.ZN (n_0_138_4), .A (sps__n55));
INV_X1 i_0_138_9 (.ZN (n_0_138_3), .A (sps__n28));
INV_X1 i_0_138_8 (.ZN (n_0_138_2), .A (sps__n43));
INV_X1 i_0_138_7 (.ZN (n_0_138_1), .A (sps__n92));
NAND4_X1 i_0_138_2 (.ZN (n_0_138_0), .A1 (n_0_138_4), .A2 (n_0_138_3), .A3 (n_0_138_2), .A4 (n_0_138_1));
NAND3_X1 i_0_121_31 (.ZN (n_0_121_30), .A1 (n_0_121_27), .A2 (n_0_121_28), .A3 (n_0_121_29));
NOR2_X1 i_0_121_30 (.ZN (n_0_121_29), .A1 (n_0_121_13), .A2 (n_0_121_23));
NOR2_X1 i_0_121_29 (.ZN (n_0_121_28), .A1 (n_0_121_22), .A2 (n_0_121_21));
NOR2_X1 i_0_121_28 (.ZN (n_0_121_27), .A1 (n_0_121_17), .A2 (n_0_121_20));
NOR2_X1 i_0_121_27 (.ZN (n_0_121_26), .A1 (n_0_121_17), .A2 (n_0_121_13));
NOR2_X1 i_0_121_26 (.ZN (n_0_121_25), .A1 (n_0_121_20), .A2 (n_0_121_21));
NOR2_X1 i_0_121_25 (.ZN (n_0_121_24), .A1 (n_0_121_22), .A2 (n_0_121_23));
NAND3_X1 i_0_121_24 (.ZN (n_0_121_23), .A1 (n_0_121_4), .A2 (n_0_121_2), .A3 (n_0_121_6));
NAND3_X1 i_0_121_23 (.ZN (n_0_121_22), .A1 (n_0_121_1), .A2 (n_0_121_3), .A3 (n_0_121_5));
NAND3_X1 i_0_121_22 (.ZN (n_0_121_21), .A1 (n_0_121_10), .A2 (n_0_121_8), .A3 (n_0_121_12));
NAND3_X1 i_0_121_21 (.ZN (n_0_121_20), .A1 (n_0_121_7), .A2 (n_0_121_9), .A3 (n_0_121_11));
NAND2_X1 i_0_121_20 (.ZN (n_0_121_19), .A1 (n_0_121_30), .A2 (\mem[5][13] ));
INV_X1 i_0_121_19 (.ZN (n_0_121_18), .A (sps__n112));
NAND4_X1 i_0_121_18 (.ZN (n_0_121_17), .A1 (n_0_121_18), .A2 (sps__n3), .A3 (sps__n121), .A4 (sps__n97));
INV_X1 i_0_121_17 (.ZN (n_0_121_16), .A (sps__n21));
INV_X1 i_0_121_16 (.ZN (n_0_121_15), .A (sps__n80));
INV_X1 i_0_121_15 (.ZN (n_0_121_14), .A (sps__n103));
NAND3_X1 i_0_121_14 (.ZN (n_0_121_13), .A1 (n_0_121_16), .A2 (n_0_121_15), .A3 (n_0_121_14));
INV_X1 i_0_121_13 (.ZN (n_0_121_12), .A (sps__n63));
INV_X1 i_0_121_12 (.ZN (n_0_121_11), .A (sps__n74));
INV_X1 i_0_121_11 (.ZN (n_0_121_10), .A (sps__n8));
INV_X1 i_0_121_10 (.ZN (n_0_121_9), .A (sps__n14));
INV_X1 i_0_121_9 (.ZN (n_0_121_8), .A (sps__n87));
INV_X1 i_0_121_8 (.ZN (n_0_121_7), .A (sps__n34));
INV_X1 i_0_121_7 (.ZN (n_0_121_6), .A (sps__n91));
INV_X1 i_0_121_6 (.ZN (n_0_121_5), .A (sps__n68));
INV_X1 i_0_121_5 (.ZN (n_0_121_4), .A (sps__n26));
INV_X1 i_0_121_4 (.ZN (n_0_121_3), .A (sps__n44));
INV_X1 i_0_121_3 (.ZN (n_0_121_2), .A (sps__n49));
INV_X1 i_0_121_2 (.ZN (n_0_121_1), .A (sps__n57));
NAND4_X1 i_0_121_1 (.ZN (n_0_121_0), .A1 (n_0_121_26), .A2 (n_0_121_25), .A3 (n_0_121_24), .A4 (data[13]));
NAND2_X1 i_0_121_0 (.ZN (n_0_46), .A1 (n_0_121_19), .A2 (n_0_121_0));
NAND3_X1 i_0_104_31 (.ZN (n_0_104_30), .A1 (n_0_104_27), .A2 (n_0_104_28), .A3 (n_0_104_29));
NOR2_X1 i_0_104_30 (.ZN (n_0_104_29), .A1 (n_0_104_13), .A2 (n_0_104_23));
NOR2_X1 i_0_104_29 (.ZN (n_0_104_28), .A1 (n_0_104_22), .A2 (n_0_104_21));
NOR2_X1 i_0_104_28 (.ZN (n_0_104_27), .A1 (n_0_104_17), .A2 (n_0_104_20));
NOR2_X1 i_0_104_27 (.ZN (n_0_104_26), .A1 (n_0_104_17), .A2 (n_0_104_13));
NOR2_X1 i_0_104_26 (.ZN (n_0_104_25), .A1 (n_0_104_20), .A2 (n_0_104_21));
NOR2_X1 i_0_104_25 (.ZN (n_0_104_24), .A1 (n_0_104_22), .A2 (n_0_104_23));
NAND3_X1 i_0_104_24 (.ZN (n_0_104_23), .A1 (n_0_104_4), .A2 (n_0_104_2), .A3 (n_0_104_6));
NAND3_X1 i_0_104_23 (.ZN (n_0_104_22), .A1 (n_0_104_1), .A2 (n_0_104_3), .A3 (n_0_104_5));
NAND3_X1 i_0_104_22 (.ZN (n_0_104_21), .A1 (n_0_104_10), .A2 (n_0_104_8), .A3 (n_0_104_12));
NAND3_X1 i_0_104_21 (.ZN (n_0_104_20), .A1 (n_0_104_7), .A2 (n_0_104_9), .A3 (n_0_104_11));
NAND2_X1 i_0_104_20 (.ZN (n_0_104_19), .A1 (n_0_104_30), .A2 (\mem[6][13] ));
INV_X1 i_0_104_19 (.ZN (n_0_104_18), .A (sps__n98));
NAND4_X1 i_0_104_18 (.ZN (n_0_104_17), .A1 (n_0_104_18), .A2 (sps__n2), .A3 (sps__n123), .A4 (sps__n114));
INV_X1 i_0_104_17 (.ZN (n_0_104_16), .A (sps__n20));
INV_X1 i_0_104_16 (.ZN (n_0_104_15), .A (sps__n81));
INV_X1 i_0_104_15 (.ZN (n_0_104_14), .A (sps__n104));
NAND3_X1 i_0_104_14 (.ZN (n_0_104_13), .A1 (n_0_104_16), .A2 (n_0_104_15), .A3 (n_0_104_14));
INV_X1 i_0_104_13 (.ZN (n_0_104_12), .A (sps__n62));
INV_X1 i_0_104_12 (.ZN (n_0_104_11), .A (sps__n74));
INV_X1 i_0_104_11 (.ZN (n_0_104_10), .A (sps__n8));
INV_X1 i_0_104_10 (.ZN (n_0_104_9), .A (sps__n15));
INV_X1 i_0_104_9 (.ZN (n_0_104_8), .A (sps__n86));
INV_X1 i_0_104_8 (.ZN (n_0_104_7), .A (sps__n36));
INV_X1 i_0_104_7 (.ZN (n_0_104_6), .A (sps__n91));
INV_X1 i_0_104_6 (.ZN (n_0_104_5), .A (sps__n68));
INV_X1 i_0_104_5 (.ZN (n_0_104_4), .A (sps__n28));
INV_X1 i_0_104_4 (.ZN (n_0_104_3), .A (sps__n42));
INV_X1 i_0_104_3 (.ZN (n_0_104_2), .A (sps__n50));
INV_X1 i_0_104_2 (.ZN (n_0_104_1), .A (sps__n55));
NAND4_X1 i_0_104_1 (.ZN (n_0_104_0), .A1 (n_0_104_26), .A2 (n_0_104_25), .A3 (n_0_104_24), .A4 (data[13]));
NAND2_X1 i_0_104_0 (.ZN (n_0_45), .A1 (n_0_104_19), .A2 (n_0_104_0));
NAND3_X1 i_0_87_27 (.ZN (n_0_87_26), .A1 (n_0_87_23), .A2 (n_0_87_24), .A3 (n_0_87_25));
NOR2_X1 i_0_87_26 (.ZN (n_0_87_25), .A1 (n_0_87_17), .A2 (n_0_87_13));
NOR2_X1 i_0_87_25 (.ZN (n_0_87_24), .A1 (n_0_87_19), .A2 (n_0_87_20));
NOR2_X1 i_0_87_24 (.ZN (n_0_87_23), .A1 (n_0_87_21), .A2 (n_0_87_22));
NAND3_X1 i_0_87_23 (.ZN (n_0_87_22), .A1 (n_0_87_4), .A2 (n_0_87_2), .A3 (n_0_87_6));
NAND3_X1 i_0_87_22 (.ZN (n_0_87_21), .A1 (n_0_87_1), .A2 (n_0_87_3), .A3 (n_0_87_5));
NAND3_X1 i_0_87_21 (.ZN (n_0_87_20), .A1 (n_0_87_10), .A2 (n_0_87_8), .A3 (n_0_87_12));
NAND3_X1 i_0_87_20 (.ZN (n_0_87_19), .A1 (n_0_87_7), .A2 (n_0_87_9), .A3 (n_0_87_11));
NAND2_X1 i_0_87_19 (.ZN (n_0_87_18), .A1 (n_0_87_26), .A2 (\mem[7][13] ));
NAND4_X1 i_0_87_18 (.ZN (n_0_87_17), .A1 (sps__n1), .A2 (sps__n121), .A3 (sps__n113), .A4 (sps__n97));
INV_X1 i_0_87_17 (.ZN (n_0_87_16), .A (sps__n21));
INV_X1 i_0_87_16 (.ZN (n_0_87_15), .A (sps__n80));
INV_X1 i_0_87_15 (.ZN (n_0_87_14), .A (sps__n103));
NAND3_X1 i_0_87_14 (.ZN (n_0_87_13), .A1 (n_0_87_16), .A2 (n_0_87_15), .A3 (n_0_87_14));
INV_X1 i_0_87_13 (.ZN (n_0_87_12), .A (sps__n61));
INV_X1 i_0_87_12 (.ZN (n_0_87_11), .A (sps__n74));
INV_X1 i_0_87_11 (.ZN (n_0_87_10), .A (sps__n7));
INV_X1 i_0_87_10 (.ZN (n_0_87_9), .A (sps__n13));
INV_X1 i_0_87_9 (.ZN (n_0_87_8), .A (sps__n87));
INV_X1 i_0_87_8 (.ZN (n_0_87_7), .A (sps__n34));
INV_X1 i_0_87_7 (.ZN (n_0_87_6), .A (sps__n91));
INV_X1 i_0_87_6 (.ZN (n_0_87_5), .A (sps__n69));
INV_X1 i_0_87_5 (.ZN (n_0_87_4), .A (sps__n27));
INV_X1 i_0_87_4 (.ZN (n_0_87_3), .A (sps__n41));
INV_X1 i_0_87_3 (.ZN (n_0_87_2), .A (sps__n49));
INV_X1 i_0_87_2 (.ZN (n_0_87_1), .A (sps__n56));
NAND4_X1 i_0_87_1 (.ZN (n_0_87_0), .A1 (n_0_87_25), .A2 (n_0_87_24), .A3 (n_0_87_23), .A4 (data[13]));
NAND2_X1 i_0_87_0 (.ZN (n_0_44), .A1 (n_0_87_18), .A2 (n_0_87_0));
NAND3_X1 i_0_70_35 (.ZN (n_0_43), .A1 (n_0_70_32), .A2 (n_0_70_33), .A3 (n_0_70_34));
NAND2_X1 i_0_70_34 (.ZN (n_0_70_34), .A1 (n_0_70_23), .A2 (\mem[8][13] ));
NAND3_X1 i_0_70_29 (.ZN (n_0_70_33), .A1 (n_0_70_26), .A2 (n_0_70_31), .A3 (n_0_70_28));
NAND2_X1 i_0_70_28 (.ZN (n_0_70_32), .A1 (n_0_70_27), .A2 (\mem[8][13] ));
NOR2_X1 i_0_70_24 (.ZN (n_0_70_31), .A1 (n_0_70_18), .A2 (n_0_70_0));
INV_X1 i_0_70_23 (.ZN (n_0_70_30), .A (n_0_70_0));
INV_X1 i_0_70_22 (.ZN (n_0_70_29), .A (n_0_70_18));
INV_X1 i_0_70_21 (.ZN (n_0_70_28), .A (n_0_70_5));
NAND3_X1 i_0_70_20 (.ZN (n_0_70_27), .A1 (n_0_70_28), .A2 (n_0_70_30), .A3 (n_0_70_9));
NOR2_X1 i_0_70_19 (.ZN (n_0_70_26), .A1 (n_0_70_14), .A2 (n_0_70_24));
INV_X1 i_0_70_18 (.ZN (n_0_70_25), .A (n_0_70_14));
NAND2_X1 i_0_70_17 (.ZN (n_0_70_24), .A1 (n_0_70_9), .A2 (data[13]));
NAND2_X1 i_0_70_16 (.ZN (n_0_70_23), .A1 (n_0_70_29), .A2 (n_0_70_25));
INV_X1 i_0_70_33 (.ZN (n_0_70_22), .A (sps__n36));
INV_X1 i_0_70_32 (.ZN (n_0_70_21), .A (sps__n8));
INV_X1 i_0_70_31 (.ZN (n_0_70_20), .A (sps__n15));
INV_X1 i_0_70_30 (.ZN (n_0_70_19), .A (sps__n50));
NAND4_X1 i_0_70_3 (.ZN (n_0_70_18), .A1 (n_0_70_22), .A2 (n_0_70_21), .A3 (n_0_70_20), .A4 (n_0_70_19));
INV_X1 i_0_70_27 (.ZN (n_0_70_17), .A (sps__n62));
INV_X1 i_0_70_26 (.ZN (n_0_70_16), .A (sps__n74));
INV_X1 i_0_70_25 (.ZN (n_0_70_15), .A (sps__n86));
NAND4_X1 i_0_70_8 (.ZN (n_0_70_14), .A1 (n_0_70_17), .A2 (n_0_70_16), .A3 (n_0_70_15), .A4 (sps__n2));
INV_X1 i_0_70_15 (.ZN (n_0_70_13), .A (sps__n121));
INV_X1 i_0_70_14 (.ZN (n_0_70_12), .A (sps__n114));
INV_X1 i_0_70_13 (.ZN (n_0_70_11), .A (sps__n97));
NAND3_X1 i_0_70_12 (.ZN (n_0_70_10), .A1 (n_0_70_13), .A2 (n_0_70_12), .A3 (n_0_70_11));
INV_X1 i_0_70_11 (.ZN (n_0_70_9), .A (n_0_70_10));
INV_X1 i_0_70_10 (.ZN (n_0_70_8), .A (sps__n68));
INV_X1 i_0_70_9 (.ZN (n_0_70_7), .A (sps__n19));
INV_X1 i_0_70_7 (.ZN (n_0_70_6), .A (sps__n81));
NAND4_X1 i_0_70_6 (.ZN (n_0_70_5), .A1 (n_0_70_8), .A2 (n_0_70_7), .A3 (n_0_70_6), .A4 (sps__n104));
INV_X1 i_0_70_5 (.ZN (n_0_70_4), .A (sps__n55));
INV_X1 i_0_70_4 (.ZN (n_0_70_3), .A (sps__n26));
INV_X1 i_0_70_2 (.ZN (n_0_70_2), .A (sps__n44));
INV_X1 i_0_70_1 (.ZN (n_0_70_1), .A (sps__n91));
NAND4_X1 i_0_70_0 (.ZN (n_0_70_0), .A1 (n_0_70_4), .A2 (n_0_70_3), .A3 (n_0_70_2), .A4 (n_0_70_1));
NOR2_X1 i_0_53_34 (.ZN (n_0_53_33), .A1 (n_0_53_19), .A2 (n_0_53_0));
INV_X1 i_0_53_33 (.ZN (n_0_53_32), .A (n_0_53_0));
INV_X1 i_0_53_28 (.ZN (n_0_53_31), .A (n_0_53_19));
NAND2_X1 i_0_53_27 (.ZN (n_0_53_30), .A1 (n_0_53_29), .A2 (\mem[9][13] ));
NAND3_X1 i_0_53_23 (.ZN (n_0_53_29), .A1 (n_0_53_5), .A2 (n_0_53_32), .A3 (n_0_53_10));
NAND3_X1 i_0_53_22 (.ZN (n_0_53_28), .A1 (n_0_53_27), .A2 (n_0_53_33), .A3 (n_0_53_14));
NOR2_X1 i_0_53_21 (.ZN (n_0_53_27), .A1 (n_0_53_6), .A2 (n_0_53_26));
NAND2_X1 i_0_53_20 (.ZN (n_0_53_26), .A1 (n_0_53_10), .A2 (data[13]));
NAND2_X1 i_0_53_19 (.ZN (n_0_53_25), .A1 (n_0_53_31), .A2 (n_0_53_14));
NAND3_X1 i_0_53_18 (.ZN (n_0_42), .A1 (n_0_53_28), .A2 (n_0_53_30), .A3 (n_0_53_24));
NAND2_X1 i_0_53_17 (.ZN (n_0_53_24), .A1 (n_0_53_25), .A2 (\mem[9][13] ));
INV_X1 i_0_53_32 (.ZN (n_0_53_23), .A (sps__n34));
INV_X1 i_0_53_31 (.ZN (n_0_53_22), .A (sps__n8));
INV_X1 i_0_53_30 (.ZN (n_0_53_21), .A (sps__n13));
INV_X1 i_0_53_29 (.ZN (n_0_53_20), .A (sps__n49));
NAND4_X1 i_0_53_3 (.ZN (n_0_53_19), .A1 (n_0_53_23), .A2 (n_0_53_22), .A3 (n_0_53_21), .A4 (n_0_53_20));
INV_X1 i_0_53_26 (.ZN (n_0_53_18), .A (sps__n61));
INV_X1 i_0_53_25 (.ZN (n_0_53_17), .A (sps__n74));
INV_X1 i_0_53_24 (.ZN (n_0_53_16), .A (sps__n87));
NAND4_X1 i_0_53_6 (.ZN (n_0_53_15), .A1 (n_0_53_18), .A2 (n_0_53_17), .A3 (n_0_53_16), .A4 (sps__n1));
INV_X1 i_0_53_16 (.ZN (n_0_53_14), .A (n_0_53_15));
INV_X1 i_0_53_15 (.ZN (n_0_53_13), .A (sps__n121));
INV_X1 i_0_53_14 (.ZN (n_0_53_12), .A (sps__n113));
NAND3_X1 i_0_53_13 (.ZN (n_0_53_11), .A1 (n_0_53_13), .A2 (n_0_53_12), .A3 (sps__n97));
INV_X1 i_0_53_12 (.ZN (n_0_53_10), .A (n_0_53_11));
INV_X1 i_0_53_11 (.ZN (n_0_53_9), .A (sps__n68));
INV_X1 i_0_53_10 (.ZN (n_0_53_8), .A (sps__n21));
INV_X1 i_0_53_9 (.ZN (n_0_53_7), .A (sps__n80));
NAND4_X1 i_0_53_8 (.ZN (n_0_53_6), .A1 (n_0_53_9), .A2 (n_0_53_8), .A3 (n_0_53_7), .A4 (sps__n103));
INV_X1 i_0_53_7 (.ZN (n_0_53_5), .A (n_0_53_6));
INV_X1 i_0_53_5 (.ZN (n_0_53_4), .A (sps__n57));
INV_X1 i_0_53_4 (.ZN (n_0_53_3), .A (sps__n27));
INV_X1 i_0_53_2 (.ZN (n_0_53_2), .A (sps__n41));
INV_X1 i_0_53_1 (.ZN (n_0_53_1), .A (sps__n91));
NAND4_X1 i_0_53_0 (.ZN (n_0_53_0), .A1 (n_0_53_4), .A2 (n_0_53_3), .A3 (n_0_53_2), .A4 (n_0_53_1));
NOR2_X1 i_0_36_34 (.ZN (n_0_36_33), .A1 (n_0_36_19), .A2 (n_0_36_0));
INV_X1 i_0_36_33 (.ZN (n_0_36_32), .A (n_0_36_0));
INV_X1 i_0_36_28 (.ZN (n_0_36_31), .A (n_0_36_19));
NAND2_X1 i_0_36_27 (.ZN (n_0_36_30), .A1 (n_0_36_29), .A2 (\mem[10][13] ));
NAND3_X1 i_0_36_23 (.ZN (n_0_36_29), .A1 (n_0_36_5), .A2 (n_0_36_32), .A3 (n_0_36_10));
NAND3_X1 i_0_36_22 (.ZN (n_0_36_28), .A1 (n_0_36_27), .A2 (n_0_36_33), .A3 (n_0_36_14));
NOR2_X1 i_0_36_21 (.ZN (n_0_36_27), .A1 (n_0_36_6), .A2 (n_0_36_26));
NAND2_X1 i_0_36_20 (.ZN (n_0_36_26), .A1 (n_0_36_10), .A2 (data[13]));
NAND2_X1 i_0_36_19 (.ZN (n_0_36_25), .A1 (n_0_36_31), .A2 (n_0_36_14));
NAND3_X1 i_0_36_18 (.ZN (n_0_41), .A1 (n_0_36_28), .A2 (n_0_36_30), .A3 (n_0_36_24));
NAND2_X1 i_0_36_17 (.ZN (n_0_36_24), .A1 (n_0_36_25), .A2 (\mem[10][13] ));
INV_X1 i_0_36_32 (.ZN (n_0_36_23), .A (sps__n34));
INV_X1 i_0_36_31 (.ZN (n_0_36_22), .A (sps__n8));
INV_X1 i_0_36_30 (.ZN (n_0_36_21), .A (sps__n15));
INV_X1 i_0_36_29 (.ZN (n_0_36_20), .A (sps__n50));
NAND4_X1 i_0_36_3 (.ZN (n_0_36_19), .A1 (n_0_36_23), .A2 (n_0_36_22), .A3 (n_0_36_21), .A4 (n_0_36_20));
INV_X1 i_0_36_26 (.ZN (n_0_36_18), .A (sps__n62));
INV_X1 i_0_36_25 (.ZN (n_0_36_17), .A (sps__n74));
INV_X1 i_0_36_24 (.ZN (n_0_36_16), .A (sps__n86));
NAND4_X1 i_0_36_6 (.ZN (n_0_36_15), .A1 (n_0_36_18), .A2 (n_0_36_17), .A3 (n_0_36_16), .A4 (sps__n3));
INV_X1 i_0_36_16 (.ZN (n_0_36_14), .A (n_0_36_15));
INV_X1 i_0_36_15 (.ZN (n_0_36_13), .A (sps__n121));
INV_X1 i_0_36_14 (.ZN (n_0_36_12), .A (sps__n99));
NAND3_X1 i_0_36_13 (.ZN (n_0_36_11), .A1 (n_0_36_13), .A2 (n_0_36_12), .A3 (sps__n112));
INV_X1 i_0_36_12 (.ZN (n_0_36_10), .A (n_0_36_11));
INV_X1 i_0_36_11 (.ZN (n_0_36_9), .A (sps__n68));
INV_X1 i_0_36_10 (.ZN (n_0_36_8), .A (sps__n19));
INV_X1 i_0_36_9 (.ZN (n_0_36_7), .A (sps__n81));
NAND4_X1 i_0_36_8 (.ZN (n_0_36_6), .A1 (n_0_36_9), .A2 (n_0_36_8), .A3 (n_0_36_7), .A4 (sps__n104));
INV_X1 i_0_36_7 (.ZN (n_0_36_5), .A (n_0_36_6));
INV_X1 i_0_36_5 (.ZN (n_0_36_4), .A (sps__n55));
INV_X1 i_0_36_4 (.ZN (n_0_36_3), .A (sps__n28));
INV_X1 i_0_36_2 (.ZN (n_0_36_2), .A (sps__n42));
INV_X1 i_0_36_1 (.ZN (n_0_36_1), .A (sps__n91));
NAND4_X1 i_0_36_0 (.ZN (n_0_36_0), .A1 (n_0_36_4), .A2 (n_0_36_3), .A3 (n_0_36_2), .A4 (n_0_36_1));
NAND3_X1 i_0_19_37 (.ZN (n_0_40), .A1 (n_0_19_34), .A2 (n_0_19_35), .A3 (n_0_19_36));
NAND2_X1 i_0_19_36 (.ZN (n_0_19_36), .A1 (n_0_19_25), .A2 (\mem[0][14] ));
NAND3_X1 i_0_19_35 (.ZN (n_0_19_35), .A1 (n_0_19_27), .A2 (n_0_19_33), .A3 (n_0_19_30));
NAND2_X1 i_0_19_34 (.ZN (n_0_19_34), .A1 (n_0_19_24), .A2 (\mem[0][14] ));
NOR2_X1 i_0_19_33 (.ZN (n_0_19_33), .A1 (n_0_19_0), .A2 (n_0_19_19));
INV_X1 i_0_19_32 (.ZN (n_0_19_32), .A (n_0_19_19));
INV_X1 i_0_19_31 (.ZN (n_0_19_31), .A (n_0_19_0));
NOR2_X1 i_0_19_30 (.ZN (n_0_19_30), .A1 (n_0_19_5), .A2 (n_0_19_15));
INV_X1 i_0_19_29 (.ZN (n_0_19_29), .A (n_0_19_15));
INV_X1 i_0_19_28 (.ZN (n_0_19_28), .A (n_0_19_5));
INV_X1 i_0_19_27 (.ZN (n_0_19_27), .A (n_0_19_26));
NAND2_X1 i_0_19_26 (.ZN (n_0_19_26), .A1 (n_0_19_10), .A2 (data[14]));
NAND2_X1 i_0_19_25 (.ZN (n_0_19_25), .A1 (n_0_19_31), .A2 (n_0_19_28));
NAND3_X1 i_0_19_24 (.ZN (n_0_19_24), .A1 (n_0_19_32), .A2 (n_0_19_29), .A3 (n_0_19_10));
INV_X1 i_0_19_23 (.ZN (n_0_19_23), .A (sps__n36));
INV_X1 i_0_19_22 (.ZN (n_0_19_22), .A (sps__n7));
INV_X1 i_0_19_21 (.ZN (n_0_19_21), .A (address[12]));
INV_X1 i_0_19_20 (.ZN (n_0_19_20), .A (sps__n49));
NAND4_X1 i_0_19_19 (.ZN (n_0_19_19), .A1 (n_0_19_23), .A2 (n_0_19_22), .A3 (n_0_19_21), .A4 (n_0_19_20));
INV_X1 i_0_19_18 (.ZN (n_0_19_18), .A (sps__n61));
INV_X1 i_0_19_17 (.ZN (n_0_19_17), .A (sps__n73));
INV_X1 i_0_19_12 (.ZN (n_0_19_16), .A (sps__n85));
NAND4_X1 i_0_19_11 (.ZN (n_0_19_15), .A1 (n_0_19_18), .A2 (n_0_19_17), .A3 (n_0_19_16), .A4 (sps__n1));
INV_X1 i_0_19_6 (.ZN (n_0_19_14), .A (address[2]));
INV_X1 i_0_19_5 (.ZN (n_0_19_13), .A (sps__n113));
INV_X1 i_0_19_4 (.ZN (n_0_19_12), .A (sps__n97));
NAND3_X1 i_0_19_1 (.ZN (n_0_19_11), .A1 (n_0_19_14), .A2 (n_0_19_13), .A3 (n_0_19_12));
INV_X1 i_0_19_0 (.ZN (n_0_19_10), .A (n_0_19_11));
INV_X1 i_0_19_16 (.ZN (n_0_19_9), .A (sps__n69));
INV_X1 i_0_19_15 (.ZN (n_0_19_8), .A (sps__n20));
INV_X1 i_0_19_14 (.ZN (n_0_19_7), .A (sps__n79));
INV_X1 i_0_19_13 (.ZN (n_0_19_6), .A (sps__n103));
NAND4_X1 i_0_19_3 (.ZN (n_0_19_5), .A1 (n_0_19_9), .A2 (n_0_19_8), .A3 (n_0_19_7), .A4 (n_0_19_6));
INV_X1 i_0_19_10 (.ZN (n_0_19_4), .A (sps__n56));
INV_X1 i_0_19_9 (.ZN (n_0_19_3), .A (sps__n27));
INV_X1 i_0_19_8 (.ZN (n_0_19_2), .A (sps__n41));
INV_X1 i_0_19_7 (.ZN (n_0_19_1), .A (sps__n93));
NAND4_X1 i_0_19_2 (.ZN (n_0_19_0), .A1 (n_0_19_4), .A2 (n_0_19_3), .A3 (n_0_19_2), .A4 (n_0_19_1));
NAND3_X1 i_0_33_36 (.ZN (n_0_39), .A1 (n_0_33_33), .A2 (n_0_33_34), .A3 (n_0_33_35));
NAND2_X1 i_0_33_35 (.ZN (n_0_33_35), .A1 (n_0_33_24), .A2 (\mem[1][14] ));
NAND2_X1 i_0_33_34 (.ZN (n_0_33_34), .A1 (n_0_33_23), .A2 (\mem[1][14] ));
NAND3_X1 i_0_33_33 (.ZN (n_0_33_33), .A1 (n_0_33_26), .A2 (n_0_33_32), .A3 (n_0_33_29));
NOR2_X1 i_0_33_32 (.ZN (n_0_33_32), .A1 (n_0_33_0), .A2 (n_0_33_18));
INV_X1 i_0_33_31 (.ZN (n_0_33_31), .A (n_0_33_18));
INV_X1 i_0_33_30 (.ZN (n_0_33_30), .A (n_0_33_0));
NOR2_X1 i_0_33_29 (.ZN (n_0_33_29), .A1 (n_0_33_5), .A2 (n_0_33_14));
INV_X1 i_0_33_28 (.ZN (n_0_33_28), .A (n_0_33_14));
INV_X1 i_0_33_27 (.ZN (n_0_33_27), .A (n_0_33_5));
INV_X1 i_0_33_26 (.ZN (n_0_33_26), .A (n_0_33_25));
NAND2_X1 i_0_33_25 (.ZN (n_0_33_25), .A1 (n_0_33_10), .A2 (data[14]));
NAND2_X1 i_0_33_24 (.ZN (n_0_33_24), .A1 (n_0_33_30), .A2 (n_0_33_27));
NAND3_X1 i_0_33_23 (.ZN (n_0_33_23), .A1 (n_0_33_31), .A2 (n_0_33_28), .A3 (n_0_33_10));
INV_X1 i_0_33_22 (.ZN (n_0_33_22), .A (sps__n35));
INV_X1 i_0_33_21 (.ZN (n_0_33_21), .A (sps__n8));
INV_X1 i_0_33_20 (.ZN (n_0_33_20), .A (sps__n13));
INV_X1 i_0_33_19 (.ZN (n_0_33_19), .A (sps__n49));
NAND4_X1 i_0_33_18 (.ZN (n_0_33_18), .A1 (n_0_33_22), .A2 (n_0_33_21), .A3 (n_0_33_20), .A4 (n_0_33_19));
INV_X1 i_0_33_17 (.ZN (n_0_33_17), .A (sps__n61));
INV_X1 i_0_33_12 (.ZN (n_0_33_16), .A (sps__n73));
INV_X1 i_0_33_11 (.ZN (n_0_33_15), .A (sps__n85));
NAND4_X1 i_0_33_6 (.ZN (n_0_33_14), .A1 (n_0_33_17), .A2 (n_0_33_16), .A3 (n_0_33_15), .A4 (sps__n1));
INV_X1 i_0_33_5 (.ZN (n_0_33_13), .A (sps__n121));
INV_X1 i_0_33_4 (.ZN (n_0_33_12), .A (sps__n112));
NAND3_X1 i_0_33_1 (.ZN (n_0_33_11), .A1 (n_0_33_13), .A2 (n_0_33_12), .A3 (sps__n97));
INV_X1 i_0_33_0 (.ZN (n_0_33_10), .A (n_0_33_11));
INV_X1 i_0_33_16 (.ZN (n_0_33_9), .A (sps__n67));
INV_X1 i_0_33_15 (.ZN (n_0_33_8), .A (sps__n21));
INV_X1 i_0_33_14 (.ZN (n_0_33_7), .A (sps__n79));
INV_X1 i_0_33_13 (.ZN (n_0_33_6), .A (sps__n106));
NAND4_X1 i_0_33_3 (.ZN (n_0_33_5), .A1 (n_0_33_9), .A2 (n_0_33_8), .A3 (n_0_33_7), .A4 (n_0_33_6));
INV_X1 i_0_33_10 (.ZN (n_0_33_4), .A (sps__n57));
INV_X1 i_0_33_9 (.ZN (n_0_33_3), .A (sps__n27));
INV_X1 i_0_33_8 (.ZN (n_0_33_2), .A (sps__n44));
INV_X1 i_0_33_7 (.ZN (n_0_33_1), .A (sps__n93));
NAND4_X1 i_0_33_2 (.ZN (n_0_33_0), .A1 (n_0_33_4), .A2 (n_0_33_3), .A3 (n_0_33_2), .A4 (n_0_33_1));
NAND3_X1 i_0_171_36 (.ZN (n_0_38), .A1 (n_0_171_33), .A2 (n_0_171_34), .A3 (n_0_171_35));
NAND2_X1 i_0_171_35 (.ZN (n_0_171_35), .A1 (n_0_171_24), .A2 (\mem[2][14] ));
NAND2_X1 i_0_171_34 (.ZN (n_0_171_34), .A1 (n_0_171_23), .A2 (\mem[2][14] ));
NAND3_X1 i_0_171_33 (.ZN (n_0_171_33), .A1 (n_0_171_26), .A2 (n_0_171_32), .A3 (n_0_171_29));
NOR2_X1 i_0_171_32 (.ZN (n_0_171_32), .A1 (n_0_171_0), .A2 (n_0_171_18));
INV_X1 i_0_171_31 (.ZN (n_0_171_31), .A (n_0_171_18));
INV_X1 i_0_171_30 (.ZN (n_0_171_30), .A (n_0_171_0));
NOR2_X1 i_0_171_29 (.ZN (n_0_171_29), .A1 (n_0_171_5), .A2 (n_0_171_14));
INV_X1 i_0_171_28 (.ZN (n_0_171_28), .A (n_0_171_14));
INV_X1 i_0_171_27 (.ZN (n_0_171_27), .A (n_0_171_5));
INV_X1 i_0_171_26 (.ZN (n_0_171_26), .A (n_0_171_25));
NAND2_X1 i_0_171_25 (.ZN (n_0_171_25), .A1 (n_0_171_10), .A2 (data[14]));
NAND2_X1 i_0_171_24 (.ZN (n_0_171_24), .A1 (n_0_171_30), .A2 (n_0_171_27));
NAND3_X1 i_0_171_23 (.ZN (n_0_171_23), .A1 (n_0_171_31), .A2 (n_0_171_28), .A3 (n_0_171_10));
INV_X1 i_0_171_22 (.ZN (n_0_171_22), .A (sps__n36));
INV_X1 i_0_171_21 (.ZN (n_0_171_21), .A (sps__n7));
INV_X1 i_0_171_20 (.ZN (n_0_171_20), .A (sps__n13));
INV_X1 i_0_171_19 (.ZN (n_0_171_19), .A (sps__n49));
NAND4_X1 i_0_171_18 (.ZN (n_0_171_18), .A1 (n_0_171_22), .A2 (n_0_171_21), .A3 (n_0_171_20), .A4 (n_0_171_19));
INV_X1 i_0_171_17 (.ZN (n_0_171_17), .A (sps__n61));
INV_X1 i_0_171_12 (.ZN (n_0_171_16), .A (sps__n73));
INV_X1 i_0_171_11 (.ZN (n_0_171_15), .A (sps__n85));
NAND4_X1 i_0_171_6 (.ZN (n_0_171_14), .A1 (n_0_171_17), .A2 (n_0_171_16), .A3 (n_0_171_15), .A4 (sps__n1));
INV_X1 i_0_171_5 (.ZN (n_0_171_13), .A (address[2]));
INV_X1 i_0_171_4 (.ZN (n_0_171_12), .A (sps__n97));
NAND3_X1 i_0_171_1 (.ZN (n_0_171_11), .A1 (n_0_171_13), .A2 (n_0_171_12), .A3 (sps__n113));
INV_X1 i_0_171_0 (.ZN (n_0_171_10), .A (n_0_171_11));
INV_X1 i_0_171_16 (.ZN (n_0_171_9), .A (sps__n69));
INV_X1 i_0_171_15 (.ZN (n_0_171_8), .A (sps__n21));
INV_X1 i_0_171_14 (.ZN (n_0_171_7), .A (sps__n79));
INV_X1 i_0_171_13 (.ZN (n_0_171_6), .A (sps__n103));
NAND4_X1 i_0_171_3 (.ZN (n_0_171_5), .A1 (n_0_171_9), .A2 (n_0_171_8), .A3 (n_0_171_7), .A4 (n_0_171_6));
INV_X1 i_0_171_10 (.ZN (n_0_171_4), .A (sps__n56));
INV_X1 i_0_171_9 (.ZN (n_0_171_3), .A (sps__n27));
INV_X1 i_0_171_8 (.ZN (n_0_171_2), .A (sps__n41));
INV_X1 i_0_171_7 (.ZN (n_0_171_1), .A (sps__n91));
NAND4_X1 i_0_171_2 (.ZN (n_0_171_0), .A1 (n_0_171_4), .A2 (n_0_171_3), .A3 (n_0_171_2), .A4 (n_0_171_1));
NAND3_X1 i_0_154_31 (.ZN (n_0_154_30), .A1 (n_0_154_27), .A2 (n_0_154_28), .A3 (n_0_154_29));
NOR2_X1 i_0_154_30 (.ZN (n_0_154_29), .A1 (n_0_154_13), .A2 (n_0_154_23));
NOR2_X1 i_0_154_29 (.ZN (n_0_154_28), .A1 (n_0_154_22), .A2 (n_0_154_21));
NOR2_X1 i_0_154_28 (.ZN (n_0_154_27), .A1 (n_0_154_17), .A2 (n_0_154_20));
NOR2_X1 i_0_154_27 (.ZN (n_0_154_26), .A1 (n_0_154_17), .A2 (n_0_154_13));
NOR2_X1 i_0_154_26 (.ZN (n_0_154_25), .A1 (n_0_154_20), .A2 (n_0_154_21));
NOR2_X1 i_0_154_25 (.ZN (n_0_154_24), .A1 (n_0_154_22), .A2 (n_0_154_23));
NAND3_X1 i_0_154_24 (.ZN (n_0_154_23), .A1 (n_0_154_4), .A2 (n_0_154_2), .A3 (n_0_154_6));
NAND3_X1 i_0_154_23 (.ZN (n_0_154_22), .A1 (n_0_154_1), .A2 (n_0_154_3), .A3 (n_0_154_5));
NAND3_X1 i_0_154_22 (.ZN (n_0_154_21), .A1 (n_0_154_10), .A2 (n_0_154_8), .A3 (n_0_154_12));
NAND3_X1 i_0_154_21 (.ZN (n_0_154_20), .A1 (n_0_154_7), .A2 (n_0_154_9), .A3 (n_0_154_11));
NAND2_X1 i_0_154_20 (.ZN (n_0_154_19), .A1 (n_0_154_30), .A2 (\mem[3][14] ));
INV_X1 i_0_154_19 (.ZN (n_0_154_18), .A (sps__n121));
NAND4_X1 i_0_154_18 (.ZN (n_0_154_17), .A1 (n_0_154_18), .A2 (sps__n1), .A3 (sps__n112), .A4 (sps__n97));
INV_X1 i_0_154_17 (.ZN (n_0_154_16), .A (sps__n21));
INV_X1 i_0_154_16 (.ZN (n_0_154_15), .A (sps__n80));
INV_X1 i_0_154_15 (.ZN (n_0_154_14), .A (sps__n103));
NAND3_X1 i_0_154_14 (.ZN (n_0_154_13), .A1 (n_0_154_16), .A2 (n_0_154_15), .A3 (n_0_154_14));
INV_X1 i_0_154_13 (.ZN (n_0_154_12), .A (sps__n61));
INV_X1 i_0_154_12 (.ZN (n_0_154_11), .A (sps__n74));
INV_X1 i_0_154_11 (.ZN (n_0_154_10), .A (sps__n8));
INV_X1 i_0_154_10 (.ZN (n_0_154_9), .A (sps__n13));
INV_X1 i_0_154_9 (.ZN (n_0_154_8), .A (sps__n87));
INV_X1 i_0_154_8 (.ZN (n_0_154_7), .A (sps__n34));
INV_X1 i_0_154_7 (.ZN (n_0_154_6), .A (sps__n93));
INV_X1 i_0_154_6 (.ZN (n_0_154_5), .A (sps__n67));
INV_X1 i_0_154_5 (.ZN (n_0_154_4), .A (sps__n27));
INV_X1 i_0_154_4 (.ZN (n_0_154_3), .A (sps__n44));
INV_X1 i_0_154_3 (.ZN (n_0_154_2), .A (sps__n49));
INV_X1 i_0_154_2 (.ZN (n_0_154_1), .A (sps__n57));
NAND4_X1 i_0_154_1 (.ZN (n_0_154_0), .A1 (n_0_154_26), .A2 (n_0_154_25), .A3 (n_0_154_24), .A4 (data[14]));
NAND2_X1 i_0_154_0 (.ZN (n_0_37), .A1 (n_0_154_19), .A2 (n_0_154_0));
NAND3_X1 i_0_137_36 (.ZN (n_0_36), .A1 (n_0_137_33), .A2 (n_0_137_34), .A3 (n_0_137_35));
NAND2_X1 i_0_137_35 (.ZN (n_0_137_35), .A1 (n_0_137_24), .A2 (\mem[4][14] ));
NAND2_X1 i_0_137_34 (.ZN (n_0_137_34), .A1 (n_0_137_23), .A2 (\mem[4][14] ));
NAND3_X1 i_0_137_33 (.ZN (n_0_137_33), .A1 (n_0_137_26), .A2 (n_0_137_32), .A3 (n_0_137_29));
NOR2_X1 i_0_137_32 (.ZN (n_0_137_32), .A1 (n_0_137_0), .A2 (n_0_137_18));
INV_X1 i_0_137_31 (.ZN (n_0_137_31), .A (n_0_137_18));
INV_X1 i_0_137_30 (.ZN (n_0_137_30), .A (n_0_137_0));
NOR2_X1 i_0_137_29 (.ZN (n_0_137_29), .A1 (n_0_137_5), .A2 (n_0_137_14));
INV_X1 i_0_137_28 (.ZN (n_0_137_28), .A (n_0_137_14));
INV_X1 i_0_137_27 (.ZN (n_0_137_27), .A (n_0_137_5));
INV_X1 i_0_137_26 (.ZN (n_0_137_26), .A (n_0_137_25));
NAND2_X1 i_0_137_25 (.ZN (n_0_137_25), .A1 (n_0_137_10), .A2 (data[14]));
NAND2_X1 i_0_137_24 (.ZN (n_0_137_24), .A1 (n_0_137_30), .A2 (n_0_137_27));
NAND3_X1 i_0_137_23 (.ZN (n_0_137_23), .A1 (n_0_137_31), .A2 (n_0_137_28), .A3 (n_0_137_10));
INV_X1 i_0_137_22 (.ZN (n_0_137_22), .A (sps__n36));
INV_X1 i_0_137_21 (.ZN (n_0_137_21), .A (sps__n7));
INV_X1 i_0_137_20 (.ZN (n_0_137_20), .A (address[12]));
INV_X1 i_0_137_19 (.ZN (n_0_137_19), .A (sps__n49));
NAND4_X1 i_0_137_18 (.ZN (n_0_137_18), .A1 (n_0_137_22), .A2 (n_0_137_21), .A3 (n_0_137_20), .A4 (n_0_137_19));
INV_X1 i_0_137_17 (.ZN (n_0_137_17), .A (sps__n61));
INV_X1 i_0_137_12 (.ZN (n_0_137_16), .A (sps__n74));
INV_X1 i_0_137_11 (.ZN (n_0_137_15), .A (sps__n87));
NAND4_X1 i_0_137_6 (.ZN (n_0_137_14), .A1 (n_0_137_17), .A2 (n_0_137_16), .A3 (n_0_137_15), .A4 (sps__n1));
INV_X1 i_0_137_5 (.ZN (n_0_137_13), .A (sps__n114));
INV_X1 i_0_137_4 (.ZN (n_0_137_12), .A (sps__n97));
NAND3_X1 i_0_137_1 (.ZN (n_0_137_11), .A1 (n_0_137_13), .A2 (n_0_137_12), .A3 (address[2]));
INV_X1 i_0_137_0 (.ZN (n_0_137_10), .A (n_0_137_11));
INV_X1 i_0_137_16 (.ZN (n_0_137_9), .A (sps__n69));
INV_X1 i_0_137_15 (.ZN (n_0_137_8), .A (sps__n20));
INV_X1 i_0_137_14 (.ZN (n_0_137_7), .A (sps__n79));
INV_X1 i_0_137_13 (.ZN (n_0_137_6), .A (sps__n103));
NAND4_X1 i_0_137_3 (.ZN (n_0_137_5), .A1 (n_0_137_9), .A2 (n_0_137_8), .A3 (n_0_137_7), .A4 (n_0_137_6));
INV_X1 i_0_137_10 (.ZN (n_0_137_4), .A (sps__n56));
INV_X1 i_0_137_9 (.ZN (n_0_137_3), .A (sps__n27));
INV_X1 i_0_137_8 (.ZN (n_0_137_2), .A (sps__n41));
INV_X1 i_0_137_7 (.ZN (n_0_137_1), .A (sps__n91));
NAND4_X1 i_0_137_2 (.ZN (n_0_137_0), .A1 (n_0_137_4), .A2 (n_0_137_3), .A3 (n_0_137_2), .A4 (n_0_137_1));
NAND3_X1 i_0_120_31 (.ZN (n_0_120_30), .A1 (n_0_120_27), .A2 (n_0_120_28), .A3 (n_0_120_29));
NOR2_X1 i_0_120_30 (.ZN (n_0_120_29), .A1 (n_0_120_13), .A2 (n_0_120_23));
NOR2_X1 i_0_120_29 (.ZN (n_0_120_28), .A1 (n_0_120_22), .A2 (n_0_120_21));
NOR2_X1 i_0_120_28 (.ZN (n_0_120_27), .A1 (n_0_120_17), .A2 (n_0_120_20));
NOR2_X1 i_0_120_27 (.ZN (n_0_120_26), .A1 (n_0_120_17), .A2 (n_0_120_13));
NOR2_X1 i_0_120_26 (.ZN (n_0_120_25), .A1 (n_0_120_20), .A2 (n_0_120_21));
NOR2_X1 i_0_120_25 (.ZN (n_0_120_24), .A1 (n_0_120_22), .A2 (n_0_120_23));
NAND3_X1 i_0_120_24 (.ZN (n_0_120_23), .A1 (n_0_120_4), .A2 (n_0_120_2), .A3 (n_0_120_6));
NAND3_X1 i_0_120_23 (.ZN (n_0_120_22), .A1 (n_0_120_1), .A2 (n_0_120_3), .A3 (n_0_120_5));
NAND3_X1 i_0_120_22 (.ZN (n_0_120_21), .A1 (n_0_120_10), .A2 (n_0_120_8), .A3 (n_0_120_12));
NAND3_X1 i_0_120_21 (.ZN (n_0_120_20), .A1 (n_0_120_7), .A2 (n_0_120_9), .A3 (n_0_120_11));
NAND2_X1 i_0_120_20 (.ZN (n_0_120_19), .A1 (n_0_120_30), .A2 (\mem[5][14] ));
INV_X1 i_0_120_19 (.ZN (n_0_120_18), .A (sps__n112));
NAND4_X1 i_0_120_18 (.ZN (n_0_120_17), .A1 (n_0_120_18), .A2 (sps__n1), .A3 (sps__n121), .A4 (sps__n97));
INV_X1 i_0_120_17 (.ZN (n_0_120_16), .A (sps__n21));
INV_X1 i_0_120_16 (.ZN (n_0_120_15), .A (sps__n80));
INV_X1 i_0_120_15 (.ZN (n_0_120_14), .A (sps__n103));
NAND3_X1 i_0_120_14 (.ZN (n_0_120_13), .A1 (n_0_120_16), .A2 (n_0_120_15), .A3 (n_0_120_14));
INV_X1 i_0_120_13 (.ZN (n_0_120_12), .A (sps__n63));
INV_X1 i_0_120_12 (.ZN (n_0_120_11), .A (sps__n74));
INV_X1 i_0_120_11 (.ZN (n_0_120_10), .A (sps__n8));
INV_X1 i_0_120_10 (.ZN (n_0_120_9), .A (sps__n13));
INV_X1 i_0_120_9 (.ZN (n_0_120_8), .A (sps__n87));
INV_X1 i_0_120_8 (.ZN (n_0_120_7), .A (sps__n35));
INV_X1 i_0_120_7 (.ZN (n_0_120_6), .A (sps__n93));
INV_X1 i_0_120_6 (.ZN (n_0_120_5), .A (sps__n67));
INV_X1 i_0_120_5 (.ZN (n_0_120_4), .A (sps__n27));
INV_X1 i_0_120_4 (.ZN (n_0_120_3), .A (sps__n44));
INV_X1 i_0_120_3 (.ZN (n_0_120_2), .A (sps__n49));
INV_X1 i_0_120_2 (.ZN (n_0_120_1), .A (sps__n57));
NAND4_X1 i_0_120_1 (.ZN (n_0_120_0), .A1 (n_0_120_26), .A2 (n_0_120_25), .A3 (n_0_120_24), .A4 (data[14]));
NAND2_X1 i_0_120_0 (.ZN (n_0_35), .A1 (n_0_120_19), .A2 (n_0_120_0));
NAND3_X1 i_0_103_31 (.ZN (n_0_103_30), .A1 (n_0_103_27), .A2 (n_0_103_28), .A3 (n_0_103_29));
NOR2_X1 i_0_103_30 (.ZN (n_0_103_29), .A1 (n_0_103_13), .A2 (n_0_103_23));
NOR2_X1 i_0_103_29 (.ZN (n_0_103_28), .A1 (n_0_103_22), .A2 (n_0_103_21));
NOR2_X1 i_0_103_28 (.ZN (n_0_103_27), .A1 (n_0_103_17), .A2 (n_0_103_20));
NOR2_X1 i_0_103_27 (.ZN (n_0_103_26), .A1 (n_0_103_17), .A2 (n_0_103_13));
NOR2_X1 i_0_103_26 (.ZN (n_0_103_25), .A1 (n_0_103_20), .A2 (n_0_103_21));
NOR2_X1 i_0_103_25 (.ZN (n_0_103_24), .A1 (n_0_103_22), .A2 (n_0_103_23));
NAND3_X1 i_0_103_24 (.ZN (n_0_103_23), .A1 (n_0_103_4), .A2 (n_0_103_2), .A3 (n_0_103_6));
NAND3_X1 i_0_103_23 (.ZN (n_0_103_22), .A1 (n_0_103_1), .A2 (n_0_103_3), .A3 (n_0_103_5));
NAND3_X1 i_0_103_22 (.ZN (n_0_103_21), .A1 (n_0_103_10), .A2 (n_0_103_8), .A3 (n_0_103_12));
NAND3_X1 i_0_103_21 (.ZN (n_0_103_20), .A1 (n_0_103_7), .A2 (n_0_103_9), .A3 (n_0_103_11));
NAND2_X1 i_0_103_20 (.ZN (n_0_103_19), .A1 (n_0_103_30), .A2 (\mem[6][14] ));
INV_X1 i_0_103_19 (.ZN (n_0_103_18), .A (sps__n97));
NAND4_X1 i_0_103_18 (.ZN (n_0_103_17), .A1 (n_0_103_18), .A2 (sps__n1), .A3 (sps__n119), .A4 (sps__n113));
INV_X1 i_0_103_17 (.ZN (n_0_103_16), .A (sps__n21));
INV_X1 i_0_103_16 (.ZN (n_0_103_15), .A (sps__n79));
INV_X1 i_0_103_15 (.ZN (n_0_103_14), .A (sps__n106));
NAND3_X1 i_0_103_14 (.ZN (n_0_103_13), .A1 (n_0_103_16), .A2 (n_0_103_15), .A3 (n_0_103_14));
INV_X1 i_0_103_13 (.ZN (n_0_103_12), .A (sps__n61));
INV_X1 i_0_103_12 (.ZN (n_0_103_11), .A (read_signal));
INV_X1 i_0_103_11 (.ZN (n_0_103_10), .A (sps__n7));
INV_X1 i_0_103_10 (.ZN (n_0_103_9), .A (sps__n13));
INV_X1 i_0_103_9 (.ZN (n_0_103_8), .A (sps__n85));
INV_X1 i_0_103_8 (.ZN (n_0_103_7), .A (sps__n36));
INV_X1 i_0_103_7 (.ZN (n_0_103_6), .A (sps__n93));
INV_X1 i_0_103_6 (.ZN (n_0_103_5), .A (sps__n69));
INV_X1 i_0_103_5 (.ZN (n_0_103_4), .A (sps__n27));
INV_X1 i_0_103_4 (.ZN (n_0_103_3), .A (sps__n41));
INV_X1 i_0_103_3 (.ZN (n_0_103_2), .A (address[11]));
INV_X1 i_0_103_2 (.ZN (n_0_103_1), .A (sps__n56));
NAND4_X1 i_0_103_1 (.ZN (n_0_103_0), .A1 (n_0_103_26), .A2 (n_0_103_25), .A3 (n_0_103_24), .A4 (data[14]));
NAND2_X1 i_0_103_0 (.ZN (n_0_34), .A1 (n_0_103_19), .A2 (n_0_103_0));
NAND3_X1 i_0_86_27 (.ZN (n_0_86_26), .A1 (n_0_86_23), .A2 (n_0_86_24), .A3 (n_0_86_25));
NOR2_X1 i_0_86_26 (.ZN (n_0_86_25), .A1 (n_0_86_17), .A2 (n_0_86_13));
NOR2_X1 i_0_86_25 (.ZN (n_0_86_24), .A1 (n_0_86_19), .A2 (n_0_86_20));
NOR2_X1 i_0_86_24 (.ZN (n_0_86_23), .A1 (n_0_86_21), .A2 (n_0_86_22));
NAND3_X1 i_0_86_23 (.ZN (n_0_86_22), .A1 (n_0_86_4), .A2 (n_0_86_2), .A3 (n_0_86_6));
NAND3_X1 i_0_86_22 (.ZN (n_0_86_21), .A1 (n_0_86_1), .A2 (n_0_86_3), .A3 (n_0_86_5));
NAND3_X1 i_0_86_21 (.ZN (n_0_86_20), .A1 (n_0_86_10), .A2 (n_0_86_8), .A3 (n_0_86_12));
NAND3_X1 i_0_86_20 (.ZN (n_0_86_19), .A1 (n_0_86_7), .A2 (n_0_86_9), .A3 (n_0_86_11));
NAND2_X1 i_0_86_19 (.ZN (n_0_86_18), .A1 (n_0_86_26), .A2 (\mem[7][14] ));
NAND4_X1 i_0_86_18 (.ZN (n_0_86_17), .A1 (sps__n1), .A2 (sps__n121), .A3 (sps__n112), .A4 (sps__n97));
INV_X1 i_0_86_17 (.ZN (n_0_86_16), .A (sps__n21));
INV_X1 i_0_86_16 (.ZN (n_0_86_15), .A (sps__n79));
INV_X1 i_0_86_15 (.ZN (n_0_86_14), .A (sps__n106));
NAND3_X1 i_0_86_14 (.ZN (n_0_86_13), .A1 (n_0_86_16), .A2 (n_0_86_15), .A3 (n_0_86_14));
INV_X1 i_0_86_13 (.ZN (n_0_86_12), .A (sps__n61));
INV_X1 i_0_86_12 (.ZN (n_0_86_11), .A (sps__n73));
INV_X1 i_0_86_11 (.ZN (n_0_86_10), .A (sps__n7));
INV_X1 i_0_86_10 (.ZN (n_0_86_9), .A (sps__n13));
INV_X1 i_0_86_9 (.ZN (n_0_86_8), .A (sps__n85));
INV_X1 i_0_86_8 (.ZN (n_0_86_7), .A (sps__n34));
INV_X1 i_0_86_7 (.ZN (n_0_86_6), .A (sps__n93));
INV_X1 i_0_86_6 (.ZN (n_0_86_5), .A (sps__n67));
INV_X1 i_0_86_5 (.ZN (n_0_86_4), .A (sps__n27));
INV_X1 i_0_86_4 (.ZN (n_0_86_3), .A (sps__n44));
INV_X1 i_0_86_3 (.ZN (n_0_86_2), .A (sps__n49));
INV_X1 i_0_86_2 (.ZN (n_0_86_1), .A (sps__n57));
NAND4_X1 i_0_86_1 (.ZN (n_0_86_0), .A1 (n_0_86_25), .A2 (n_0_86_24), .A3 (n_0_86_23), .A4 (data[14]));
NAND2_X1 i_0_86_0 (.ZN (n_0_33), .A1 (n_0_86_18), .A2 (n_0_86_0));
NAND3_X1 i_0_69_35 (.ZN (n_0_30), .A1 (n_0_69_32), .A2 (n_0_69_33), .A3 (n_0_69_34));
NAND2_X1 i_0_69_34 (.ZN (n_0_69_34), .A1 (n_0_69_23), .A2 (\mem[8][14] ));
NAND3_X1 i_0_69_29 (.ZN (n_0_69_33), .A1 (n_0_69_26), .A2 (n_0_69_31), .A3 (n_0_69_28));
NAND2_X1 i_0_69_28 (.ZN (n_0_69_32), .A1 (n_0_69_27), .A2 (\mem[8][14] ));
NOR2_X1 i_0_69_24 (.ZN (n_0_69_31), .A1 (n_0_69_18), .A2 (n_0_69_0));
INV_X1 i_0_69_23 (.ZN (n_0_69_30), .A (n_0_69_0));
INV_X1 i_0_69_22 (.ZN (n_0_69_29), .A (n_0_69_18));
INV_X1 i_0_69_21 (.ZN (n_0_69_28), .A (n_0_69_5));
NAND3_X1 i_0_69_20 (.ZN (n_0_69_27), .A1 (n_0_69_28), .A2 (n_0_69_30), .A3 (n_0_69_9));
NOR2_X1 i_0_69_19 (.ZN (n_0_69_26), .A1 (n_0_69_14), .A2 (n_0_69_24));
INV_X1 i_0_69_18 (.ZN (n_0_69_25), .A (n_0_69_14));
NAND2_X1 i_0_69_17 (.ZN (n_0_69_24), .A1 (n_0_69_9), .A2 (data[14]));
NAND2_X1 i_0_69_16 (.ZN (n_0_69_23), .A1 (n_0_69_29), .A2 (n_0_69_25));
INV_X1 i_0_69_33 (.ZN (n_0_69_22), .A (sps__n36));
INV_X1 i_0_69_32 (.ZN (n_0_69_21), .A (sps__n7));
INV_X1 i_0_69_31 (.ZN (n_0_69_20), .A (sps__n13));
INV_X1 i_0_69_30 (.ZN (n_0_69_19), .A (address[11]));
NAND4_X1 i_0_69_3 (.ZN (n_0_69_18), .A1 (n_0_69_22), .A2 (n_0_69_21), .A3 (n_0_69_20), .A4 (n_0_69_19));
INV_X1 i_0_69_27 (.ZN (n_0_69_17), .A (sps__n61));
INV_X1 i_0_69_26 (.ZN (n_0_69_16), .A (read_signal));
INV_X1 i_0_69_25 (.ZN (n_0_69_15), .A (address[15]));
NAND4_X1 i_0_69_8 (.ZN (n_0_69_14), .A1 (n_0_69_17), .A2 (n_0_69_16), .A3 (n_0_69_15), .A4 (write_signal));
INV_X1 i_0_69_15 (.ZN (n_0_69_13), .A (address[2]));
INV_X1 i_0_69_14 (.ZN (n_0_69_12), .A (sps__n113));
INV_X1 i_0_69_13 (.ZN (n_0_69_11), .A (address[0]));
NAND3_X1 i_0_69_12 (.ZN (n_0_69_10), .A1 (n_0_69_13), .A2 (n_0_69_12), .A3 (n_0_69_11));
INV_X1 i_0_69_11 (.ZN (n_0_69_9), .A (n_0_69_10));
INV_X1 i_0_69_10 (.ZN (n_0_69_8), .A (sps__n69));
INV_X1 i_0_69_9 (.ZN (n_0_69_7), .A (sps__n21));
INV_X1 i_0_69_7 (.ZN (n_0_69_6), .A (sps__n79));
NAND4_X1 i_0_69_6 (.ZN (n_0_69_5), .A1 (n_0_69_8), .A2 (n_0_69_7), .A3 (n_0_69_6), .A4 (sps__n106));
INV_X1 i_0_69_5 (.ZN (n_0_69_4), .A (sps__n56));
INV_X1 i_0_69_4 (.ZN (n_0_69_3), .A (sps__n27));
INV_X1 i_0_69_2 (.ZN (n_0_69_2), .A (sps__n41));
INV_X1 i_0_69_1 (.ZN (n_0_69_1), .A (sps__n93));
NAND4_X1 i_0_69_0 (.ZN (n_0_69_0), .A1 (n_0_69_4), .A2 (n_0_69_3), .A3 (n_0_69_2), .A4 (n_0_69_1));
NOR2_X1 i_0_52_34 (.ZN (n_0_52_33), .A1 (n_0_52_19), .A2 (n_0_52_0));
INV_X1 i_0_52_33 (.ZN (n_0_52_32), .A (n_0_52_0));
INV_X1 i_0_52_28 (.ZN (n_0_52_31), .A (n_0_52_19));
NAND2_X1 i_0_52_27 (.ZN (n_0_52_30), .A1 (n_0_52_29), .A2 (\mem[9][14] ));
NAND3_X1 i_0_52_23 (.ZN (n_0_52_29), .A1 (n_0_52_5), .A2 (n_0_52_32), .A3 (n_0_52_10));
NAND3_X1 i_0_52_22 (.ZN (n_0_52_28), .A1 (n_0_52_27), .A2 (n_0_52_33), .A3 (n_0_52_14));
NOR2_X1 i_0_52_21 (.ZN (n_0_52_27), .A1 (n_0_52_6), .A2 (n_0_52_26));
NAND2_X1 i_0_52_20 (.ZN (n_0_52_26), .A1 (n_0_52_10), .A2 (data[14]));
NAND2_X1 i_0_52_19 (.ZN (n_0_52_25), .A1 (n_0_52_31), .A2 (n_0_52_14));
NAND3_X1 i_0_52_18 (.ZN (n_0_29), .A1 (n_0_52_28), .A2 (n_0_52_30), .A3 (n_0_52_24));
NAND2_X1 i_0_52_17 (.ZN (n_0_52_24), .A1 (n_0_52_25), .A2 (\mem[9][14] ));
INV_X1 i_0_52_32 (.ZN (n_0_52_23), .A (sps__n34));
INV_X1 i_0_52_31 (.ZN (n_0_52_22), .A (sps__n7));
INV_X1 i_0_52_30 (.ZN (n_0_52_21), .A (sps__n13));
INV_X1 i_0_52_29 (.ZN (n_0_52_20), .A (sps__n49));
NAND4_X1 i_0_52_3 (.ZN (n_0_52_19), .A1 (n_0_52_23), .A2 (n_0_52_22), .A3 (n_0_52_21), .A4 (n_0_52_20));
INV_X1 i_0_52_26 (.ZN (n_0_52_18), .A (sps__n61));
INV_X1 i_0_52_25 (.ZN (n_0_52_17), .A (sps__n73));
INV_X1 i_0_52_24 (.ZN (n_0_52_16), .A (sps__n85));
NAND4_X1 i_0_52_6 (.ZN (n_0_52_15), .A1 (n_0_52_18), .A2 (n_0_52_17), .A3 (n_0_52_16), .A4 (sps__n1));
INV_X1 i_0_52_16 (.ZN (n_0_52_14), .A (n_0_52_15));
INV_X1 i_0_52_15 (.ZN (n_0_52_13), .A (sps__n119));
INV_X1 i_0_52_14 (.ZN (n_0_52_12), .A (sps__n113));
NAND3_X1 i_0_52_13 (.ZN (n_0_52_11), .A1 (n_0_52_13), .A2 (n_0_52_12), .A3 (sps__n97));
INV_X1 i_0_52_12 (.ZN (n_0_52_10), .A (n_0_52_11));
INV_X1 i_0_52_11 (.ZN (n_0_52_9), .A (sps__n67));
INV_X1 i_0_52_10 (.ZN (n_0_52_8), .A (sps__n21));
INV_X1 i_0_52_9 (.ZN (n_0_52_7), .A (sps__n79));
NAND4_X1 i_0_52_8 (.ZN (n_0_52_6), .A1 (n_0_52_9), .A2 (n_0_52_8), .A3 (n_0_52_7), .A4 (sps__n106));
INV_X1 i_0_52_7 (.ZN (n_0_52_5), .A (n_0_52_6));
INV_X1 i_0_52_5 (.ZN (n_0_52_4), .A (sps__n56));
INV_X1 i_0_52_4 (.ZN (n_0_52_3), .A (sps__n27));
INV_X1 i_0_52_2 (.ZN (n_0_52_2), .A (sps__n41));
INV_X1 i_0_52_1 (.ZN (n_0_52_1), .A (sps__n93));
NAND4_X1 i_0_52_0 (.ZN (n_0_52_0), .A1 (n_0_52_4), .A2 (n_0_52_3), .A3 (n_0_52_2), .A4 (n_0_52_1));
NOR2_X1 i_0_35_34 (.ZN (n_0_35_33), .A1 (n_0_35_19), .A2 (n_0_35_0));
INV_X1 i_0_35_33 (.ZN (n_0_35_32), .A (n_0_35_0));
INV_X1 i_0_35_28 (.ZN (n_0_35_31), .A (n_0_35_19));
NAND2_X1 i_0_35_27 (.ZN (n_0_35_30), .A1 (n_0_35_29), .A2 (\mem[10][14] ));
NAND3_X1 i_0_35_23 (.ZN (n_0_35_29), .A1 (n_0_35_5), .A2 (n_0_35_32), .A3 (n_0_35_10));
NAND3_X1 i_0_35_22 (.ZN (n_0_35_28), .A1 (n_0_35_27), .A2 (n_0_35_33), .A3 (n_0_35_14));
NOR2_X1 i_0_35_21 (.ZN (n_0_35_27), .A1 (n_0_35_6), .A2 (n_0_35_26));
NAND2_X1 i_0_35_20 (.ZN (n_0_35_26), .A1 (n_0_35_10), .A2 (data[14]));
NAND2_X1 i_0_35_19 (.ZN (n_0_35_25), .A1 (n_0_35_31), .A2 (n_0_35_14));
NAND3_X1 i_0_35_18 (.ZN (n_0_28), .A1 (n_0_35_28), .A2 (n_0_35_30), .A3 (n_0_35_24));
NAND2_X1 i_0_35_17 (.ZN (n_0_35_24), .A1 (n_0_35_25), .A2 (\mem[10][14] ));
INV_X1 i_0_35_32 (.ZN (n_0_35_23), .A (sps__n36));
INV_X1 i_0_35_31 (.ZN (n_0_35_22), .A (sps__n7));
INV_X1 i_0_35_30 (.ZN (n_0_35_21), .A (sps__n13));
INV_X1 i_0_35_29 (.ZN (n_0_35_20), .A (sps__n49));
NAND4_X1 i_0_35_3 (.ZN (n_0_35_19), .A1 (n_0_35_23), .A2 (n_0_35_22), .A3 (n_0_35_21), .A4 (n_0_35_20));
INV_X1 i_0_35_26 (.ZN (n_0_35_18), .A (sps__n61));
INV_X1 i_0_35_25 (.ZN (n_0_35_17), .A (sps__n73));
INV_X1 i_0_35_24 (.ZN (n_0_35_16), .A (sps__n85));
NAND4_X1 i_0_35_6 (.ZN (n_0_35_15), .A1 (n_0_35_18), .A2 (n_0_35_17), .A3 (n_0_35_16), .A4 (sps__n1));
INV_X1 i_0_35_16 (.ZN (n_0_35_14), .A (n_0_35_15));
INV_X1 i_0_35_15 (.ZN (n_0_35_13), .A (address[2]));
INV_X1 i_0_35_14 (.ZN (n_0_35_12), .A (sps__n97));
NAND3_X1 i_0_35_13 (.ZN (n_0_35_11), .A1 (n_0_35_13), .A2 (n_0_35_12), .A3 (sps__n113));
INV_X1 i_0_35_12 (.ZN (n_0_35_10), .A (n_0_35_11));
INV_X1 i_0_35_11 (.ZN (n_0_35_9), .A (sps__n69));
INV_X1 i_0_35_10 (.ZN (n_0_35_8), .A (sps__n21));
INV_X1 i_0_35_9 (.ZN (n_0_35_7), .A (sps__n79));
NAND4_X1 i_0_35_8 (.ZN (n_0_35_6), .A1 (n_0_35_9), .A2 (n_0_35_8), .A3 (n_0_35_7), .A4 (sps__n103));
INV_X1 i_0_35_7 (.ZN (n_0_35_5), .A (n_0_35_6));
INV_X1 i_0_35_5 (.ZN (n_0_35_4), .A (sps__n56));
INV_X1 i_0_35_4 (.ZN (n_0_35_3), .A (sps__n27));
INV_X1 i_0_35_2 (.ZN (n_0_35_2), .A (sps__n41));
INV_X1 i_0_35_1 (.ZN (n_0_35_1), .A (sps__n93));
NAND4_X1 i_0_35_0 (.ZN (n_0_35_0), .A1 (n_0_35_4), .A2 (n_0_35_3), .A3 (n_0_35_2), .A4 (n_0_35_1));
NAND3_X1 i_0_18_37 (.ZN (n_0_27), .A1 (n_0_18_34), .A2 (n_0_18_35), .A3 (n_0_18_36));
NAND2_X1 i_0_18_36 (.ZN (n_0_18_36), .A1 (n_0_18_25), .A2 (\mem[0][15] ));
NAND3_X1 i_0_18_35 (.ZN (n_0_18_35), .A1 (n_0_18_27), .A2 (n_0_18_33), .A3 (n_0_18_30));
NAND2_X1 i_0_18_34 (.ZN (n_0_18_34), .A1 (n_0_18_24), .A2 (\mem[0][15] ));
NOR2_X1 i_0_18_33 (.ZN (n_0_18_33), .A1 (n_0_18_0), .A2 (n_0_18_19));
INV_X1 i_0_18_32 (.ZN (n_0_18_32), .A (n_0_18_19));
INV_X1 i_0_18_31 (.ZN (n_0_18_31), .A (n_0_18_0));
NOR2_X1 i_0_18_30 (.ZN (n_0_18_30), .A1 (n_0_18_5), .A2 (n_0_18_15));
INV_X1 i_0_18_29 (.ZN (n_0_18_29), .A (n_0_18_15));
INV_X1 i_0_18_28 (.ZN (n_0_18_28), .A (n_0_18_5));
INV_X1 i_0_18_27 (.ZN (n_0_18_27), .A (n_0_18_26));
NAND2_X1 i_0_18_26 (.ZN (n_0_18_26), .A1 (n_0_18_10), .A2 (data[15]));
NAND2_X1 i_0_18_25 (.ZN (n_0_18_25), .A1 (n_0_18_31), .A2 (n_0_18_28));
NAND3_X1 i_0_18_24 (.ZN (n_0_18_24), .A1 (n_0_18_32), .A2 (n_0_18_29), .A3 (n_0_18_10));
INV_X1 i_0_18_23 (.ZN (n_0_18_23), .A (sps__n36));
INV_X1 i_0_18_22 (.ZN (n_0_18_22), .A (sps__n7));
INV_X1 i_0_18_21 (.ZN (n_0_18_21), .A (sps__n14));
INV_X1 i_0_18_20 (.ZN (n_0_18_20), .A (sps__n49));
NAND4_X1 i_0_18_19 (.ZN (n_0_18_19), .A1 (n_0_18_23), .A2 (n_0_18_22), .A3 (n_0_18_21), .A4 (n_0_18_20));
INV_X1 i_0_18_18 (.ZN (n_0_18_18), .A (RST));
INV_X1 i_0_18_17 (.ZN (n_0_18_17), .A (sps__n73));
INV_X1 i_0_18_12 (.ZN (n_0_18_16), .A (sps__n85));
NAND4_X1 i_0_18_11 (.ZN (n_0_18_15), .A1 (n_0_18_18), .A2 (n_0_18_17), .A3 (n_0_18_16), .A4 (sps__n2));
INV_X1 i_0_18_6 (.ZN (n_0_18_14), .A (sps__n123));
INV_X1 i_0_18_5 (.ZN (n_0_18_13), .A (sps__n114));
INV_X1 i_0_18_4 (.ZN (n_0_18_12), .A (sps__n98));
NAND3_X1 i_0_18_1 (.ZN (n_0_18_11), .A1 (n_0_18_14), .A2 (n_0_18_13), .A3 (n_0_18_12));
INV_X1 i_0_18_0 (.ZN (n_0_18_10), .A (n_0_18_11));
INV_X1 i_0_18_16 (.ZN (n_0_18_9), .A (sps__n69));
INV_X1 i_0_18_15 (.ZN (n_0_18_8), .A (sps__n20));
INV_X1 i_0_18_14 (.ZN (n_0_18_7), .A (sps__n79));
INV_X1 i_0_18_13 (.ZN (n_0_18_6), .A (address[3]));
NAND4_X1 i_0_18_3 (.ZN (n_0_18_5), .A1 (n_0_18_9), .A2 (n_0_18_8), .A3 (n_0_18_7), .A4 (n_0_18_6));
INV_X1 i_0_18_10 (.ZN (n_0_18_4), .A (sps__n56));
INV_X1 i_0_18_9 (.ZN (n_0_18_3), .A (sps__n26));
INV_X1 i_0_18_8 (.ZN (n_0_18_2), .A (address[8]));
INV_X1 i_0_18_7 (.ZN (n_0_18_1), .A (address[7]));
NAND4_X1 i_0_18_2 (.ZN (n_0_18_0), .A1 (n_0_18_4), .A2 (n_0_18_3), .A3 (n_0_18_2), .A4 (n_0_18_1));
NAND3_X1 i_0_170_36 (.ZN (n_0_26), .A1 (n_0_170_33), .A2 (n_0_170_34), .A3 (n_0_170_35));
NAND2_X1 i_0_170_35 (.ZN (n_0_170_35), .A1 (n_0_170_24), .A2 (\mem[1][15] ));
NAND2_X1 i_0_170_34 (.ZN (n_0_170_34), .A1 (n_0_170_23), .A2 (\mem[1][15] ));
NAND3_X1 i_0_170_33 (.ZN (n_0_170_33), .A1 (n_0_170_26), .A2 (n_0_170_32), .A3 (n_0_170_29));
NOR2_X1 i_0_170_32 (.ZN (n_0_170_32), .A1 (n_0_170_0), .A2 (n_0_170_18));
INV_X1 i_0_170_31 (.ZN (n_0_170_31), .A (n_0_170_18));
INV_X1 i_0_170_30 (.ZN (n_0_170_30), .A (n_0_170_0));
NOR2_X1 i_0_170_29 (.ZN (n_0_170_29), .A1 (n_0_170_5), .A2 (n_0_170_14));
INV_X1 i_0_170_28 (.ZN (n_0_170_28), .A (n_0_170_14));
INV_X1 i_0_170_27 (.ZN (n_0_170_27), .A (n_0_170_5));
INV_X1 i_0_170_26 (.ZN (n_0_170_26), .A (n_0_170_25));
NAND2_X1 i_0_170_25 (.ZN (n_0_170_25), .A1 (n_0_170_10), .A2 (data[15]));
NAND2_X1 i_0_170_24 (.ZN (n_0_170_24), .A1 (n_0_170_30), .A2 (n_0_170_27));
NAND3_X1 i_0_170_23 (.ZN (n_0_170_23), .A1 (n_0_170_31), .A2 (n_0_170_28), .A3 (n_0_170_10));
INV_X1 i_0_170_22 (.ZN (n_0_170_22), .A (sps__n36));
INV_X1 i_0_170_21 (.ZN (n_0_170_21), .A (sps__n7));
INV_X1 i_0_170_20 (.ZN (n_0_170_20), .A (address[12]));
INV_X1 i_0_170_19 (.ZN (n_0_170_19), .A (sps__n49));
NAND4_X1 i_0_170_18 (.ZN (n_0_170_18), .A1 (n_0_170_22), .A2 (n_0_170_21), .A3 (n_0_170_20), .A4 (n_0_170_19));
INV_X1 i_0_170_17 (.ZN (n_0_170_17), .A (RST));
INV_X1 i_0_170_12 (.ZN (n_0_170_16), .A (sps__n73));
INV_X1 i_0_170_11 (.ZN (n_0_170_15), .A (sps__n85));
NAND4_X1 i_0_170_6 (.ZN (n_0_170_14), .A1 (n_0_170_17), .A2 (n_0_170_16), .A3 (n_0_170_15), .A4 (sps__n1));
INV_X1 i_0_170_5 (.ZN (n_0_170_13), .A (sps__n123));
INV_X1 i_0_170_4 (.ZN (n_0_170_12), .A (sps__n114));
NAND3_X1 i_0_170_1 (.ZN (n_0_170_11), .A1 (n_0_170_13), .A2 (n_0_170_12), .A3 (sps__n97));
INV_X1 i_0_170_0 (.ZN (n_0_170_10), .A (n_0_170_11));
INV_X1 i_0_170_16 (.ZN (n_0_170_9), .A (sps__n69));
INV_X1 i_0_170_15 (.ZN (n_0_170_8), .A (sps__n20));
INV_X1 i_0_170_14 (.ZN (n_0_170_7), .A (sps__n79));
INV_X1 i_0_170_13 (.ZN (n_0_170_6), .A (address[3]));
NAND4_X1 i_0_170_3 (.ZN (n_0_170_5), .A1 (n_0_170_9), .A2 (n_0_170_8), .A3 (n_0_170_7), .A4 (n_0_170_6));
INV_X1 i_0_170_10 (.ZN (n_0_170_4), .A (sps__n56));
INV_X1 i_0_170_9 (.ZN (n_0_170_3), .A (sps__n26));
INV_X1 i_0_170_8 (.ZN (n_0_170_2), .A (address[8]));
INV_X1 i_0_170_7 (.ZN (n_0_170_1), .A (address[7]));
NAND4_X1 i_0_170_2 (.ZN (n_0_170_0), .A1 (n_0_170_4), .A2 (n_0_170_3), .A3 (n_0_170_2), .A4 (n_0_170_1));
NAND3_X1 i_0_153_36 (.ZN (n_0_25), .A1 (n_0_153_33), .A2 (n_0_153_34), .A3 (n_0_153_35));
NAND2_X1 i_0_153_35 (.ZN (n_0_153_35), .A1 (n_0_153_24), .A2 (\mem[2][15] ));
NAND2_X1 i_0_153_34 (.ZN (n_0_153_34), .A1 (n_0_153_23), .A2 (\mem[2][15] ));
NAND3_X1 i_0_153_33 (.ZN (n_0_153_33), .A1 (n_0_153_26), .A2 (n_0_153_32), .A3 (n_0_153_29));
NOR2_X1 i_0_153_32 (.ZN (n_0_153_32), .A1 (n_0_153_0), .A2 (n_0_153_18));
INV_X1 i_0_153_31 (.ZN (n_0_153_31), .A (n_0_153_18));
INV_X1 i_0_153_30 (.ZN (n_0_153_30), .A (n_0_153_0));
NOR2_X1 i_0_153_29 (.ZN (n_0_153_29), .A1 (n_0_153_5), .A2 (n_0_153_14));
INV_X1 i_0_153_28 (.ZN (n_0_153_28), .A (n_0_153_14));
INV_X1 i_0_153_27 (.ZN (n_0_153_27), .A (n_0_153_5));
INV_X1 i_0_153_26 (.ZN (n_0_153_26), .A (n_0_153_25));
NAND2_X1 i_0_153_25 (.ZN (n_0_153_25), .A1 (n_0_153_10), .A2 (data[15]));
NAND2_X1 i_0_153_24 (.ZN (n_0_153_24), .A1 (n_0_153_30), .A2 (n_0_153_27));
NAND3_X1 i_0_153_23 (.ZN (n_0_153_23), .A1 (n_0_153_31), .A2 (n_0_153_28), .A3 (n_0_153_10));
INV_X1 i_0_153_22 (.ZN (n_0_153_22), .A (sps__n36));
INV_X1 i_0_153_21 (.ZN (n_0_153_21), .A (sps__n7));
INV_X1 i_0_153_20 (.ZN (n_0_153_20), .A (sps__n14));
INV_X1 i_0_153_19 (.ZN (n_0_153_19), .A (sps__n50));
NAND4_X1 i_0_153_18 (.ZN (n_0_153_18), .A1 (n_0_153_22), .A2 (n_0_153_21), .A3 (n_0_153_20), .A4 (n_0_153_19));
INV_X1 i_0_153_17 (.ZN (n_0_153_17), .A (RST));
INV_X1 i_0_153_12 (.ZN (n_0_153_16), .A (sps__n73));
INV_X1 i_0_153_11 (.ZN (n_0_153_15), .A (sps__n85));
NAND4_X1 i_0_153_6 (.ZN (n_0_153_14), .A1 (n_0_153_17), .A2 (n_0_153_16), .A3 (n_0_153_15), .A4 (sps__n2));
INV_X1 i_0_153_5 (.ZN (n_0_153_13), .A (sps__n123));
INV_X1 i_0_153_4 (.ZN (n_0_153_12), .A (sps__n98));
NAND3_X1 i_0_153_1 (.ZN (n_0_153_11), .A1 (n_0_153_13), .A2 (n_0_153_12), .A3 (sps__n114));
INV_X1 i_0_153_0 (.ZN (n_0_153_10), .A (n_0_153_11));
INV_X1 i_0_153_16 (.ZN (n_0_153_9), .A (sps__n69));
INV_X1 i_0_153_15 (.ZN (n_0_153_8), .A (sps__n20));
INV_X1 i_0_153_14 (.ZN (n_0_153_7), .A (sps__n79));
INV_X1 i_0_153_13 (.ZN (n_0_153_6), .A (address[3]));
NAND4_X1 i_0_153_3 (.ZN (n_0_153_5), .A1 (n_0_153_9), .A2 (n_0_153_8), .A3 (n_0_153_7), .A4 (n_0_153_6));
INV_X1 i_0_153_10 (.ZN (n_0_153_4), .A (sps__n56));
INV_X1 i_0_153_9 (.ZN (n_0_153_3), .A (sps__n26));
INV_X1 i_0_153_8 (.ZN (n_0_153_2), .A (address[8]));
INV_X1 i_0_153_7 (.ZN (n_0_153_1), .A (address[7]));
NAND4_X1 i_0_153_2 (.ZN (n_0_153_0), .A1 (n_0_153_4), .A2 (n_0_153_3), .A3 (n_0_153_2), .A4 (n_0_153_1));
NAND3_X1 i_0_136_31 (.ZN (n_0_136_30), .A1 (n_0_136_27), .A2 (n_0_136_28), .A3 (n_0_136_29));
NOR2_X1 i_0_136_30 (.ZN (n_0_136_29), .A1 (n_0_136_13), .A2 (n_0_136_23));
NOR2_X1 i_0_136_29 (.ZN (n_0_136_28), .A1 (n_0_136_22), .A2 (n_0_136_21));
NOR2_X1 i_0_136_28 (.ZN (n_0_136_27), .A1 (n_0_136_17), .A2 (n_0_136_20));
NOR2_X1 i_0_136_27 (.ZN (n_0_136_26), .A1 (n_0_136_17), .A2 (n_0_136_13));
NOR2_X1 i_0_136_26 (.ZN (n_0_136_25), .A1 (n_0_136_20), .A2 (n_0_136_21));
NOR2_X1 i_0_136_25 (.ZN (n_0_136_24), .A1 (n_0_136_22), .A2 (n_0_136_23));
NAND3_X1 i_0_136_24 (.ZN (n_0_136_23), .A1 (n_0_136_4), .A2 (n_0_136_2), .A3 (n_0_136_6));
NAND3_X1 i_0_136_23 (.ZN (n_0_136_22), .A1 (n_0_136_1), .A2 (n_0_136_3), .A3 (n_0_136_5));
NAND3_X1 i_0_136_22 (.ZN (n_0_136_21), .A1 (n_0_136_10), .A2 (n_0_136_8), .A3 (n_0_136_12));
NAND3_X1 i_0_136_21 (.ZN (n_0_136_20), .A1 (n_0_136_7), .A2 (n_0_136_9), .A3 (n_0_136_11));
NAND2_X1 i_0_136_20 (.ZN (n_0_136_19), .A1 (n_0_136_30), .A2 (\mem[3][15] ));
INV_X1 i_0_136_19 (.ZN (n_0_136_18), .A (sps__n123));
NAND4_X1 i_0_136_18 (.ZN (n_0_136_17), .A1 (n_0_136_18), .A2 (sps__n2), .A3 (sps__n114), .A4 (sps__n98));
INV_X1 i_0_136_17 (.ZN (n_0_136_16), .A (sps__n20));
INV_X1 i_0_136_16 (.ZN (n_0_136_15), .A (sps__n80));
INV_X1 i_0_136_15 (.ZN (n_0_136_14), .A (sps__n103));
NAND3_X1 i_0_136_14 (.ZN (n_0_136_13), .A1 (n_0_136_16), .A2 (n_0_136_15), .A3 (n_0_136_14));
INV_X1 i_0_136_13 (.ZN (n_0_136_12), .A (sps__n61));
INV_X1 i_0_136_12 (.ZN (n_0_136_11), .A (sps__n74));
INV_X1 i_0_136_11 (.ZN (n_0_136_10), .A (sps__n7));
INV_X1 i_0_136_10 (.ZN (n_0_136_9), .A (sps__n14));
INV_X1 i_0_136_9 (.ZN (n_0_136_8), .A (sps__n85));
INV_X1 i_0_136_8 (.ZN (n_0_136_7), .A (sps__n36));
INV_X1 i_0_136_7 (.ZN (n_0_136_6), .A (sps__n91));
INV_X1 i_0_136_6 (.ZN (n_0_136_5), .A (sps__n69));
INV_X1 i_0_136_5 (.ZN (n_0_136_4), .A (sps__n26));
INV_X1 i_0_136_4 (.ZN (n_0_136_3), .A (sps__n44));
INV_X1 i_0_136_3 (.ZN (n_0_136_2), .A (sps__n50));
INV_X1 i_0_136_2 (.ZN (n_0_136_1), .A (sps__n56));
NAND4_X1 i_0_136_1 (.ZN (n_0_136_0), .A1 (n_0_136_26), .A2 (n_0_136_25), .A3 (n_0_136_24), .A4 (data[15]));
NAND2_X1 i_0_136_0 (.ZN (n_0_24), .A1 (n_0_136_19), .A2 (n_0_136_0));
NAND3_X1 i_0_119_36 (.ZN (n_0_23), .A1 (n_0_119_33), .A2 (n_0_119_34), .A3 (n_0_119_35));
NAND2_X1 i_0_119_35 (.ZN (n_0_119_35), .A1 (n_0_119_24), .A2 (\mem[4][15] ));
NAND2_X1 i_0_119_34 (.ZN (n_0_119_34), .A1 (n_0_119_23), .A2 (\mem[4][15] ));
NAND3_X1 i_0_119_33 (.ZN (n_0_119_33), .A1 (n_0_119_26), .A2 (n_0_119_32), .A3 (n_0_119_29));
NOR2_X1 i_0_119_32 (.ZN (n_0_119_32), .A1 (n_0_119_0), .A2 (n_0_119_18));
INV_X1 i_0_119_31 (.ZN (n_0_119_31), .A (n_0_119_18));
INV_X1 i_0_119_30 (.ZN (n_0_119_30), .A (n_0_119_0));
NOR2_X1 i_0_119_29 (.ZN (n_0_119_29), .A1 (n_0_119_5), .A2 (n_0_119_14));
INV_X1 i_0_119_28 (.ZN (n_0_119_28), .A (n_0_119_14));
INV_X1 i_0_119_27 (.ZN (n_0_119_27), .A (n_0_119_5));
INV_X1 i_0_119_26 (.ZN (n_0_119_26), .A (n_0_119_25));
NAND2_X1 i_0_119_25 (.ZN (n_0_119_25), .A1 (n_0_119_10), .A2 (data[15]));
NAND2_X1 i_0_119_24 (.ZN (n_0_119_24), .A1 (n_0_119_30), .A2 (n_0_119_27));
NAND3_X1 i_0_119_23 (.ZN (n_0_119_23), .A1 (n_0_119_31), .A2 (n_0_119_28), .A3 (n_0_119_10));
INV_X1 i_0_119_22 (.ZN (n_0_119_22), .A (sps__n36));
INV_X1 i_0_119_21 (.ZN (n_0_119_21), .A (sps__n7));
INV_X1 i_0_119_20 (.ZN (n_0_119_20), .A (sps__n14));
INV_X1 i_0_119_19 (.ZN (n_0_119_19), .A (sps__n50));
NAND4_X1 i_0_119_18 (.ZN (n_0_119_18), .A1 (n_0_119_22), .A2 (n_0_119_21), .A3 (n_0_119_20), .A4 (n_0_119_19));
INV_X1 i_0_119_17 (.ZN (n_0_119_17), .A (RST));
INV_X1 i_0_119_12 (.ZN (n_0_119_16), .A (sps__n74));
INV_X1 i_0_119_11 (.ZN (n_0_119_15), .A (sps__n85));
NAND4_X1 i_0_119_6 (.ZN (n_0_119_14), .A1 (n_0_119_17), .A2 (n_0_119_16), .A3 (n_0_119_15), .A4 (sps__n2));
INV_X1 i_0_119_5 (.ZN (n_0_119_13), .A (sps__n114));
INV_X1 i_0_119_4 (.ZN (n_0_119_12), .A (sps__n98));
NAND3_X1 i_0_119_1 (.ZN (n_0_119_11), .A1 (n_0_119_13), .A2 (n_0_119_12), .A3 (sps__n123));
INV_X1 i_0_119_0 (.ZN (n_0_119_10), .A (n_0_119_11));
INV_X1 i_0_119_16 (.ZN (n_0_119_9), .A (sps__n69));
INV_X1 i_0_119_15 (.ZN (n_0_119_8), .A (sps__n20));
INV_X1 i_0_119_14 (.ZN (n_0_119_7), .A (sps__n79));
INV_X1 i_0_119_13 (.ZN (n_0_119_6), .A (sps__n103));
NAND4_X1 i_0_119_3 (.ZN (n_0_119_5), .A1 (n_0_119_9), .A2 (n_0_119_8), .A3 (n_0_119_7), .A4 (n_0_119_6));
INV_X1 i_0_119_10 (.ZN (n_0_119_4), .A (sps__n56));
INV_X1 i_0_119_9 (.ZN (n_0_119_3), .A (sps__n26));
INV_X1 i_0_119_8 (.ZN (n_0_119_2), .A (sps__n42));
INV_X1 i_0_119_7 (.ZN (n_0_119_1), .A (address[7]));
NAND4_X1 i_0_119_2 (.ZN (n_0_119_0), .A1 (n_0_119_4), .A2 (n_0_119_3), .A3 (n_0_119_2), .A4 (n_0_119_1));
NAND3_X1 i_0_102_31 (.ZN (n_0_102_30), .A1 (n_0_102_27), .A2 (n_0_102_28), .A3 (n_0_102_29));
NOR2_X1 i_0_102_30 (.ZN (n_0_102_29), .A1 (n_0_102_13), .A2 (n_0_102_23));
NOR2_X1 i_0_102_29 (.ZN (n_0_102_28), .A1 (n_0_102_22), .A2 (n_0_102_21));
NOR2_X1 i_0_102_28 (.ZN (n_0_102_27), .A1 (n_0_102_17), .A2 (n_0_102_20));
NOR2_X1 i_0_102_27 (.ZN (n_0_102_26), .A1 (n_0_102_17), .A2 (n_0_102_13));
NOR2_X1 i_0_102_26 (.ZN (n_0_102_25), .A1 (n_0_102_20), .A2 (n_0_102_21));
NOR2_X1 i_0_102_25 (.ZN (n_0_102_24), .A1 (n_0_102_22), .A2 (n_0_102_23));
NAND3_X1 i_0_102_24 (.ZN (n_0_102_23), .A1 (n_0_102_4), .A2 (n_0_102_2), .A3 (n_0_102_6));
NAND3_X1 i_0_102_23 (.ZN (n_0_102_22), .A1 (n_0_102_1), .A2 (n_0_102_3), .A3 (n_0_102_5));
NAND3_X1 i_0_102_22 (.ZN (n_0_102_21), .A1 (n_0_102_10), .A2 (n_0_102_8), .A3 (n_0_102_12));
NAND3_X1 i_0_102_21 (.ZN (n_0_102_20), .A1 (n_0_102_7), .A2 (n_0_102_9), .A3 (n_0_102_11));
NAND2_X1 i_0_102_20 (.ZN (n_0_102_19), .A1 (n_0_102_30), .A2 (\mem[5][15] ));
INV_X1 i_0_102_19 (.ZN (n_0_102_18), .A (sps__n114));
NAND4_X1 i_0_102_18 (.ZN (n_0_102_17), .A1 (n_0_102_18), .A2 (sps__n2), .A3 (sps__n123), .A4 (sps__n98));
INV_X1 i_0_102_17 (.ZN (n_0_102_16), .A (sps__n20));
INV_X1 i_0_102_16 (.ZN (n_0_102_15), .A (sps__n79));
INV_X1 i_0_102_15 (.ZN (n_0_102_14), .A (address[3]));
NAND3_X1 i_0_102_14 (.ZN (n_0_102_13), .A1 (n_0_102_16), .A2 (n_0_102_15), .A3 (n_0_102_14));
INV_X1 i_0_102_13 (.ZN (n_0_102_12), .A (RST));
INV_X1 i_0_102_12 (.ZN (n_0_102_11), .A (sps__n73));
INV_X1 i_0_102_11 (.ZN (n_0_102_10), .A (sps__n7));
INV_X1 i_0_102_10 (.ZN (n_0_102_9), .A (sps__n14));
INV_X1 i_0_102_9 (.ZN (n_0_102_8), .A (sps__n85));
INV_X1 i_0_102_8 (.ZN (n_0_102_7), .A (sps__n36));
INV_X1 i_0_102_7 (.ZN (n_0_102_6), .A (address[7]));
INV_X1 i_0_102_6 (.ZN (n_0_102_5), .A (sps__n69));
INV_X1 i_0_102_5 (.ZN (n_0_102_4), .A (sps__n26));
INV_X1 i_0_102_4 (.ZN (n_0_102_3), .A (address[8]));
INV_X1 i_0_102_3 (.ZN (n_0_102_2), .A (sps__n49));
INV_X1 i_0_102_2 (.ZN (n_0_102_1), .A (sps__n56));
NAND4_X1 i_0_102_1 (.ZN (n_0_102_0), .A1 (n_0_102_26), .A2 (n_0_102_25), .A3 (n_0_102_24), .A4 (data[15]));
NAND2_X1 i_0_102_0 (.ZN (n_0_22), .A1 (n_0_102_19), .A2 (n_0_102_0));
NAND3_X1 i_0_85_31 (.ZN (n_0_85_30), .A1 (n_0_85_27), .A2 (n_0_85_28), .A3 (n_0_85_29));
NOR2_X1 i_0_85_30 (.ZN (n_0_85_29), .A1 (n_0_85_13), .A2 (n_0_85_23));
NOR2_X1 i_0_85_29 (.ZN (n_0_85_28), .A1 (n_0_85_22), .A2 (n_0_85_21));
NOR2_X1 i_0_85_28 (.ZN (n_0_85_27), .A1 (n_0_85_17), .A2 (n_0_85_20));
NOR2_X1 i_0_85_27 (.ZN (n_0_85_26), .A1 (n_0_85_17), .A2 (n_0_85_13));
NOR2_X1 i_0_85_26 (.ZN (n_0_85_25), .A1 (n_0_85_20), .A2 (n_0_85_21));
NOR2_X1 i_0_85_25 (.ZN (n_0_85_24), .A1 (n_0_85_22), .A2 (n_0_85_23));
NAND3_X1 i_0_85_24 (.ZN (n_0_85_23), .A1 (n_0_85_4), .A2 (n_0_85_2), .A3 (n_0_85_6));
NAND3_X1 i_0_85_23 (.ZN (n_0_85_22), .A1 (n_0_85_1), .A2 (n_0_85_3), .A3 (n_0_85_5));
NAND3_X1 i_0_85_22 (.ZN (n_0_85_21), .A1 (n_0_85_10), .A2 (n_0_85_8), .A3 (n_0_85_12));
NAND3_X1 i_0_85_21 (.ZN (n_0_85_20), .A1 (n_0_85_7), .A2 (n_0_85_9), .A3 (n_0_85_11));
NAND2_X1 i_0_85_20 (.ZN (n_0_85_19), .A1 (n_0_85_30), .A2 (\mem[6][15] ));
INV_X1 i_0_85_19 (.ZN (n_0_85_18), .A (sps__n97));
NAND4_X1 i_0_85_18 (.ZN (n_0_85_17), .A1 (n_0_85_18), .A2 (sps__n1), .A3 (sps__n123), .A4 (sps__n114));
INV_X1 i_0_85_17 (.ZN (n_0_85_16), .A (sps__n20));
INV_X1 i_0_85_16 (.ZN (n_0_85_15), .A (sps__n79));
INV_X1 i_0_85_15 (.ZN (n_0_85_14), .A (sps__n103));
NAND3_X1 i_0_85_14 (.ZN (n_0_85_13), .A1 (n_0_85_16), .A2 (n_0_85_15), .A3 (n_0_85_14));
INV_X1 i_0_85_13 (.ZN (n_0_85_12), .A (sps__n61));
INV_X1 i_0_85_12 (.ZN (n_0_85_11), .A (sps__n73));
INV_X1 i_0_85_11 (.ZN (n_0_85_10), .A (sps__n7));
INV_X1 i_0_85_10 (.ZN (n_0_85_9), .A (address[12]));
INV_X1 i_0_85_9 (.ZN (n_0_85_8), .A (sps__n85));
INV_X1 i_0_85_8 (.ZN (n_0_85_7), .A (sps__n36));
INV_X1 i_0_85_7 (.ZN (n_0_85_6), .A (sps__n91));
INV_X1 i_0_85_6 (.ZN (n_0_85_5), .A (sps__n69));
INV_X1 i_0_85_5 (.ZN (n_0_85_4), .A (sps__n27));
INV_X1 i_0_85_4 (.ZN (n_0_85_3), .A (sps__n41));
INV_X1 i_0_85_3 (.ZN (n_0_85_2), .A (sps__n49));
INV_X1 i_0_85_2 (.ZN (n_0_85_1), .A (sps__n56));
NAND4_X1 i_0_85_1 (.ZN (n_0_85_0), .A1 (n_0_85_26), .A2 (n_0_85_25), .A3 (n_0_85_24), .A4 (data[15]));
NAND2_X1 i_0_85_0 (.ZN (n_0_21), .A1 (n_0_85_19), .A2 (n_0_85_0));
NAND3_X1 i_0_68_27 (.ZN (n_0_68_26), .A1 (n_0_68_23), .A2 (n_0_68_24), .A3 (n_0_68_25));
NOR2_X1 i_0_68_26 (.ZN (n_0_68_25), .A1 (n_0_68_17), .A2 (n_0_68_13));
NOR2_X1 i_0_68_25 (.ZN (n_0_68_24), .A1 (n_0_68_19), .A2 (n_0_68_20));
NOR2_X1 i_0_68_24 (.ZN (n_0_68_23), .A1 (n_0_68_21), .A2 (n_0_68_22));
NAND3_X1 i_0_68_23 (.ZN (n_0_68_22), .A1 (n_0_68_4), .A2 (n_0_68_2), .A3 (n_0_68_6));
NAND3_X1 i_0_68_22 (.ZN (n_0_68_21), .A1 (n_0_68_1), .A2 (n_0_68_3), .A3 (n_0_68_5));
NAND3_X1 i_0_68_21 (.ZN (n_0_68_20), .A1 (n_0_68_10), .A2 (n_0_68_8), .A3 (n_0_68_12));
NAND3_X1 i_0_68_20 (.ZN (n_0_68_19), .A1 (n_0_68_7), .A2 (n_0_68_9), .A3 (n_0_68_11));
NAND2_X1 i_0_68_19 (.ZN (n_0_68_18), .A1 (n_0_68_26), .A2 (\mem[7][15] ));
NAND4_X1 i_0_68_18 (.ZN (n_0_68_17), .A1 (sps__n2), .A2 (sps__n123), .A3 (sps__n114), .A4 (sps__n98));
INV_X1 i_0_68_17 (.ZN (n_0_68_16), .A (sps__n20));
INV_X1 i_0_68_16 (.ZN (n_0_68_15), .A (sps__n79));
INV_X1 i_0_68_15 (.ZN (n_0_68_14), .A (sps__n103));
NAND3_X1 i_0_68_14 (.ZN (n_0_68_13), .A1 (n_0_68_16), .A2 (n_0_68_15), .A3 (n_0_68_14));
INV_X1 i_0_68_13 (.ZN (n_0_68_12), .A (sps__n61));
INV_X1 i_0_68_12 (.ZN (n_0_68_11), .A (sps__n73));
INV_X1 i_0_68_11 (.ZN (n_0_68_10), .A (sps__n7));
INV_X1 i_0_68_10 (.ZN (n_0_68_9), .A (address[12]));
INV_X1 i_0_68_9 (.ZN (n_0_68_8), .A (sps__n85));
INV_X1 i_0_68_8 (.ZN (n_0_68_7), .A (sps__n36));
INV_X1 i_0_68_7 (.ZN (n_0_68_6), .A (address[7]));
INV_X1 i_0_68_6 (.ZN (n_0_68_5), .A (sps__n69));
INV_X1 i_0_68_5 (.ZN (n_0_68_4), .A (sps__n27));
INV_X1 i_0_68_4 (.ZN (n_0_68_3), .A (address[8]));
INV_X1 i_0_68_3 (.ZN (n_0_68_2), .A (sps__n49));
INV_X1 i_0_68_2 (.ZN (n_0_68_1), .A (sps__n56));
NAND4_X1 i_0_68_1 (.ZN (n_0_68_0), .A1 (n_0_68_25), .A2 (n_0_68_24), .A3 (n_0_68_23), .A4 (data[15]));
NAND2_X1 i_0_68_0 (.ZN (n_0_20), .A1 (n_0_68_18), .A2 (n_0_68_0));
NAND3_X1 i_0_51_35 (.ZN (n_0_19), .A1 (n_0_51_32), .A2 (n_0_51_33), .A3 (n_0_51_34));
NAND2_X1 i_0_51_34 (.ZN (n_0_51_34), .A1 (n_0_51_23), .A2 (\mem[8][15] ));
NAND3_X1 i_0_51_29 (.ZN (n_0_51_33), .A1 (n_0_51_26), .A2 (n_0_51_31), .A3 (n_0_51_28));
NAND2_X1 i_0_51_28 (.ZN (n_0_51_32), .A1 (n_0_51_27), .A2 (\mem[8][15] ));
NOR2_X1 i_0_51_24 (.ZN (n_0_51_31), .A1 (n_0_51_18), .A2 (n_0_51_0));
INV_X1 i_0_51_23 (.ZN (n_0_51_30), .A (n_0_51_0));
INV_X1 i_0_51_22 (.ZN (n_0_51_29), .A (n_0_51_18));
INV_X1 i_0_51_21 (.ZN (n_0_51_28), .A (n_0_51_5));
NAND3_X1 i_0_51_20 (.ZN (n_0_51_27), .A1 (n_0_51_28), .A2 (n_0_51_30), .A3 (n_0_51_9));
NOR2_X1 i_0_51_19 (.ZN (n_0_51_26), .A1 (n_0_51_14), .A2 (n_0_51_24));
INV_X1 i_0_51_18 (.ZN (n_0_51_25), .A (n_0_51_14));
NAND2_X1 i_0_51_17 (.ZN (n_0_51_24), .A1 (n_0_51_9), .A2 (data[15]));
NAND2_X1 i_0_51_16 (.ZN (n_0_51_23), .A1 (n_0_51_29), .A2 (n_0_51_25));
INV_X1 i_0_51_33 (.ZN (n_0_51_22), .A (sps__n36));
INV_X1 i_0_51_32 (.ZN (n_0_51_21), .A (sps__n7));
INV_X1 i_0_51_31 (.ZN (n_0_51_20), .A (sps__n14));
INV_X1 i_0_51_30 (.ZN (n_0_51_19), .A (sps__n50));
NAND4_X1 i_0_51_3 (.ZN (n_0_51_18), .A1 (n_0_51_22), .A2 (n_0_51_21), .A3 (n_0_51_20), .A4 (n_0_51_19));
INV_X1 i_0_51_27 (.ZN (n_0_51_17), .A (RST));
INV_X1 i_0_51_26 (.ZN (n_0_51_16), .A (sps__n74));
INV_X1 i_0_51_25 (.ZN (n_0_51_15), .A (sps__n85));
NAND4_X1 i_0_51_8 (.ZN (n_0_51_14), .A1 (n_0_51_17), .A2 (n_0_51_16), .A3 (n_0_51_15), .A4 (sps__n2));
INV_X1 i_0_51_15 (.ZN (n_0_51_13), .A (sps__n123));
INV_X1 i_0_51_14 (.ZN (n_0_51_12), .A (sps__n114));
INV_X1 i_0_51_13 (.ZN (n_0_51_11), .A (sps__n98));
NAND3_X1 i_0_51_12 (.ZN (n_0_51_10), .A1 (n_0_51_13), .A2 (n_0_51_12), .A3 (n_0_51_11));
INV_X1 i_0_51_11 (.ZN (n_0_51_9), .A (n_0_51_10));
INV_X1 i_0_51_10 (.ZN (n_0_51_8), .A (sps__n69));
INV_X1 i_0_51_9 (.ZN (n_0_51_7), .A (sps__n20));
INV_X1 i_0_51_7 (.ZN (n_0_51_6), .A (sps__n80));
NAND4_X1 i_0_51_6 (.ZN (n_0_51_5), .A1 (n_0_51_8), .A2 (n_0_51_7), .A3 (n_0_51_6), .A4 (sps__n103));
INV_X1 i_0_51_5 (.ZN (n_0_51_4), .A (sps__n56));
INV_X1 i_0_51_4 (.ZN (n_0_51_3), .A (sps__n26));
INV_X1 i_0_51_2 (.ZN (n_0_51_2), .A (sps__n42));
INV_X1 i_0_51_1 (.ZN (n_0_51_1), .A (address[7]));
NAND4_X1 i_0_51_0 (.ZN (n_0_51_0), .A1 (n_0_51_4), .A2 (n_0_51_3), .A3 (n_0_51_2), .A4 (n_0_51_1));
NOR2_X1 i_0_34_34 (.ZN (n_0_34_33), .A1 (n_0_34_19), .A2 (n_0_34_0));
INV_X1 i_0_34_33 (.ZN (n_0_34_32), .A (n_0_34_0));
INV_X1 i_0_34_28 (.ZN (n_0_34_31), .A (n_0_34_19));
NAND2_X1 i_0_34_27 (.ZN (n_0_34_30), .A1 (n_0_34_29), .A2 (\mem[9][15] ));
NAND3_X1 i_0_34_23 (.ZN (n_0_34_29), .A1 (n_0_34_5), .A2 (n_0_34_32), .A3 (n_0_34_10));
NAND3_X1 i_0_34_22 (.ZN (n_0_34_28), .A1 (n_0_34_27), .A2 (n_0_34_33), .A3 (n_0_34_14));
NOR2_X1 i_0_34_21 (.ZN (n_0_34_27), .A1 (n_0_34_6), .A2 (n_0_34_26));
NAND2_X1 i_0_34_20 (.ZN (n_0_34_26), .A1 (n_0_34_10), .A2 (data[15]));
NAND2_X1 i_0_34_19 (.ZN (n_0_34_25), .A1 (n_0_34_31), .A2 (n_0_34_14));
NAND3_X1 i_0_34_18 (.ZN (n_0_18), .A1 (n_0_34_28), .A2 (n_0_34_30), .A3 (n_0_34_24));
NAND2_X1 i_0_34_17 (.ZN (n_0_34_24), .A1 (n_0_34_25), .A2 (\mem[9][15] ));
INV_X1 i_0_34_32 (.ZN (n_0_34_23), .A (sps__n36));
INV_X1 i_0_34_31 (.ZN (n_0_34_22), .A (sps__n7));
INV_X1 i_0_34_30 (.ZN (n_0_34_21), .A (sps__n14));
INV_X1 i_0_34_29 (.ZN (n_0_34_20), .A (sps__n50));
NAND4_X1 i_0_34_3 (.ZN (n_0_34_19), .A1 (n_0_34_23), .A2 (n_0_34_22), .A3 (n_0_34_21), .A4 (n_0_34_20));
INV_X1 i_0_34_26 (.ZN (n_0_34_18), .A (RST));
INV_X1 i_0_34_25 (.ZN (n_0_34_17), .A (sps__n74));
INV_X1 i_0_34_24 (.ZN (n_0_34_16), .A (sps__n85));
NAND4_X1 i_0_34_6 (.ZN (n_0_34_15), .A1 (n_0_34_18), .A2 (n_0_34_17), .A3 (n_0_34_16), .A4 (sps__n2));
INV_X1 i_0_34_16 (.ZN (n_0_34_14), .A (n_0_34_15));
INV_X1 i_0_34_15 (.ZN (n_0_34_13), .A (sps__n123));
INV_X1 i_0_34_14 (.ZN (n_0_34_12), .A (sps__n114));
NAND3_X1 i_0_34_13 (.ZN (n_0_34_11), .A1 (n_0_34_13), .A2 (n_0_34_12), .A3 (sps__n98));
INV_X1 i_0_34_12 (.ZN (n_0_34_10), .A (n_0_34_11));
INV_X1 i_0_34_11 (.ZN (n_0_34_9), .A (sps__n69));
INV_X1 i_0_34_10 (.ZN (n_0_34_8), .A (sps__n20));
INV_X1 i_0_34_9 (.ZN (n_0_34_7), .A (sps__n80));
NAND4_X1 i_0_34_8 (.ZN (n_0_34_6), .A1 (n_0_34_9), .A2 (n_0_34_8), .A3 (n_0_34_7), .A4 (sps__n103));
INV_X1 i_0_34_7 (.ZN (n_0_34_5), .A (n_0_34_6));
INV_X1 i_0_34_5 (.ZN (n_0_34_4), .A (sps__n56));
INV_X1 i_0_34_4 (.ZN (n_0_34_3), .A (sps__n26));
INV_X1 i_0_34_2 (.ZN (n_0_34_2), .A (sps__n42));
INV_X1 i_0_34_1 (.ZN (n_0_34_1), .A (sps__n91));
NAND4_X1 i_0_34_0 (.ZN (n_0_34_0), .A1 (n_0_34_4), .A2 (n_0_34_3), .A3 (n_0_34_2), .A4 (n_0_34_1));
NOR2_X1 i_0_17_34 (.ZN (n_0_17_33), .A1 (n_0_17_19), .A2 (n_0_17_0));
INV_X1 i_0_17_33 (.ZN (n_0_17_32), .A (n_0_17_0));
INV_X1 i_0_17_28 (.ZN (n_0_17_31), .A (n_0_17_19));
NAND2_X1 i_0_17_27 (.ZN (n_0_17_30), .A1 (n_0_17_29), .A2 (\mem[10][15] ));
NAND3_X1 i_0_17_23 (.ZN (n_0_17_29), .A1 (n_0_17_5), .A2 (n_0_17_32), .A3 (n_0_17_10));
NAND3_X1 i_0_17_22 (.ZN (n_0_17_28), .A1 (n_0_17_27), .A2 (n_0_17_33), .A3 (n_0_17_14));
NOR2_X1 i_0_17_21 (.ZN (n_0_17_27), .A1 (n_0_17_6), .A2 (n_0_17_26));
NAND2_X1 i_0_17_20 (.ZN (n_0_17_26), .A1 (n_0_17_10), .A2 (data[15]));
NAND2_X1 i_0_17_19 (.ZN (n_0_17_25), .A1 (n_0_17_31), .A2 (n_0_17_14));
NAND3_X1 i_0_17_18 (.ZN (n_0_17), .A1 (n_0_17_28), .A2 (n_0_17_30), .A3 (n_0_17_24));
NAND2_X1 i_0_17_17 (.ZN (n_0_17_24), .A1 (n_0_17_25), .A2 (\mem[10][15] ));
INV_X1 i_0_17_32 (.ZN (n_0_17_23), .A (sps__n36));
INV_X1 i_0_17_31 (.ZN (n_0_17_22), .A (sps__n7));
INV_X1 i_0_17_30 (.ZN (n_0_17_21), .A (address[12]));
INV_X1 i_0_17_29 (.ZN (n_0_17_20), .A (sps__n49));
NAND4_X1 i_0_17_3 (.ZN (n_0_17_19), .A1 (n_0_17_23), .A2 (n_0_17_22), .A3 (n_0_17_21), .A4 (n_0_17_20));
INV_X1 i_0_17_26 (.ZN (n_0_17_18), .A (sps__n61));
INV_X1 i_0_17_25 (.ZN (n_0_17_17), .A (sps__n74));
INV_X1 i_0_17_24 (.ZN (n_0_17_16), .A (sps__n85));
NAND4_X1 i_0_17_6 (.ZN (n_0_17_15), .A1 (n_0_17_18), .A2 (n_0_17_17), .A3 (n_0_17_16), .A4 (sps__n1));
INV_X1 i_0_17_16 (.ZN (n_0_17_14), .A (n_0_17_15));
INV_X1 i_0_17_15 (.ZN (n_0_17_13), .A (sps__n123));
INV_X1 i_0_17_14 (.ZN (n_0_17_12), .A (sps__n97));
NAND3_X1 i_0_17_13 (.ZN (n_0_17_11), .A1 (n_0_17_13), .A2 (n_0_17_12), .A3 (sps__n114));
INV_X1 i_0_17_12 (.ZN (n_0_17_10), .A (n_0_17_11));
INV_X1 i_0_17_11 (.ZN (n_0_17_9), .A (sps__n69));
INV_X1 i_0_17_10 (.ZN (n_0_17_8), .A (sps__n21));
INV_X1 i_0_17_9 (.ZN (n_0_17_7), .A (sps__n80));
NAND4_X1 i_0_17_8 (.ZN (n_0_17_6), .A1 (n_0_17_9), .A2 (n_0_17_8), .A3 (n_0_17_7), .A4 (sps__n103));
INV_X1 i_0_17_7 (.ZN (n_0_17_5), .A (n_0_17_6));
INV_X1 i_0_17_5 (.ZN (n_0_17_4), .A (sps__n56));
INV_X1 i_0_17_4 (.ZN (n_0_17_3), .A (sps__n27));
INV_X1 i_0_17_2 (.ZN (n_0_17_2), .A (sps__n41));
INV_X1 i_0_17_1 (.ZN (n_0_17_1), .A (sps__n91));
NAND4_X1 i_0_17_0 (.ZN (n_0_17_0), .A1 (n_0_17_4), .A2 (n_0_17_3), .A3 (n_0_17_2), .A4 (n_0_17_1));
INV_X1 i_0_10_35 (.ZN (n_0_10_34), .A (sps__n103));
INV_X1 i_0_10_34 (.ZN (n_0_10_33), .A (\mem[3][5] ));
INV_X1 i_0_10_33 (.ZN (n_0_10_32), .A (sps__n123));
NAND2_X1 i_0_10_32 (.ZN (n_0_10_31), .A1 (n_0_10_32), .A2 (n_0_10_33));
INV_X1 i_0_10_31 (.ZN (n_0_10_30), .A (\mem[7][5] ));
NAND2_X1 i_0_10_30 (.ZN (n_0_10_29), .A1 (sps__n123), .A2 (n_0_10_30));
NAND3_X1 i_0_10_29 (.ZN (n_0_10_28), .A1 (n_0_10_31), .A2 (n_0_10_34), .A3 (n_0_10_29));
NAND2_X1 i_0_10_28 (.ZN (n_0_10_27), .A1 (n_0_10_28), .A2 (sps__n112));
INV_X1 i_0_10_27 (.ZN (n_0_10_26), .A (sps__n112));
INV_X1 i_0_10_26 (.ZN (n_0_10_25), .A (\mem[1][5] ));
NAND2_X1 i_0_10_25 (.ZN (n_0_10_24), .A1 (n_0_10_34), .A2 (n_0_10_25));
INV_X1 i_0_10_24 (.ZN (n_0_10_23), .A (\mem[9][5] ));
NAND2_X1 i_0_10_23 (.ZN (n_0_10_22), .A1 (sps__n103), .A2 (n_0_10_23));
NAND3_X1 i_0_10_22 (.ZN (n_0_10_21), .A1 (n_0_10_24), .A2 (n_0_10_32), .A3 (n_0_10_22));
NAND3_X1 i_0_10_21 (.ZN (n_0_10_20), .A1 (n_0_10_34), .A2 (\mem[5][5] ), .A3 (sps__n123));
NAND3_X1 i_0_10_20 (.ZN (n_0_10_19), .A1 (n_0_10_21), .A2 (n_0_10_26), .A3 (n_0_10_20));
NAND3_X1 i_0_10_19 (.ZN (n_0_10_18), .A1 (n_0_10_19), .A2 (sps__n98), .A3 (n_0_10_27));
INV_X1 i_0_10_18 (.ZN (n_0_10_17), .A (sps__n98));
INV_X1 i_0_10_17 (.ZN (n_0_10_16), .A (\mem[8][5] ));
NAND2_X1 i_0_10_16 (.ZN (n_0_10_15), .A1 (n_0_10_26), .A2 (n_0_10_16));
INV_X1 i_0_10_15 (.ZN (n_0_10_14), .A (\mem[10][5] ));
NAND2_X1 i_0_10_14 (.ZN (n_0_10_13), .A1 (sps__n112), .A2 (n_0_10_14));
NAND3_X1 i_0_10_13 (.ZN (n_0_10_12), .A1 (n_0_10_15), .A2 (n_0_10_32), .A3 (n_0_10_13));
NAND2_X1 i_0_10_12 (.ZN (n_0_10_11), .A1 (n_0_10_12), .A2 (sps__n105));
NAND2_X1 i_0_10_11 (.ZN (n_0_10_10), .A1 (n_0_10_26), .A2 (\mem[0][5] ));
NAND2_X1 i_0_10_10 (.ZN (n_0_10_9), .A1 (sps__n112), .A2 (\mem[2][5] ));
NAND4_X1 i_0_10_9 (.ZN (n_0_10_8), .A1 (n_0_10_10), .A2 (n_0_10_9), .A3 (n_0_10_34), .A4 (n_0_10_32));
NAND2_X1 i_0_10_8 (.ZN (n_0_10_7), .A1 (n_0_10_26), .A2 (\mem[4][5] ));
NAND2_X1 i_0_10_7 (.ZN (n_0_10_6), .A1 (sps__n112), .A2 (\mem[6][5] ));
NAND3_X1 i_0_10_6 (.ZN (n_0_10_5), .A1 (n_0_10_7), .A2 (sps__n123), .A3 (n_0_10_6));
NAND4_X1 i_0_10_5 (.ZN (n_0_10_4), .A1 (n_0_10_11), .A2 (n_0_10_17), .A3 (n_0_10_8), .A4 (n_0_10_5));
NAND2_X1 i_0_10_4 (.ZN (n_0_10_3), .A1 (n_0_10_4), .A2 (n_0_10_18));
NAND2_X1 i_0_10_3 (.ZN (n_0_10_2), .A1 (n_0_10_3), .A2 (n_0_5));
INV_X1 i_0_10_2 (.ZN (n_0_10_1), .A (n_0_5));
NAND2_X1 i_0_10_1 (.ZN (n_0_10_0), .A1 (n_0_10_1), .A2 (dataout[5]));
NAND2_X1 i_0_10_0 (.ZN (n_0_16), .A1 (n_0_10_2), .A2 (n_0_10_0));
INV_X1 i_0_9_35 (.ZN (n_0_9_34), .A (sps__n106));
INV_X1 i_0_9_34 (.ZN (n_0_9_33), .A (\mem[3][6] ));
INV_X1 i_0_9_33 (.ZN (n_0_9_32), .A (address[2]));
NAND2_X1 i_0_9_32 (.ZN (n_0_9_31), .A1 (n_0_9_32), .A2 (n_0_9_33));
INV_X1 i_0_9_31 (.ZN (n_0_9_30), .A (\mem[7][6] ));
NAND2_X1 i_0_9_30 (.ZN (n_0_9_29), .A1 (address[2]), .A2 (n_0_9_30));
NAND3_X1 i_0_9_29 (.ZN (n_0_9_28), .A1 (n_0_9_31), .A2 (n_0_9_34), .A3 (n_0_9_29));
NAND2_X1 i_0_9_28 (.ZN (n_0_9_27), .A1 (n_0_9_28), .A2 (sps__n114));
INV_X1 i_0_9_27 (.ZN (n_0_9_26), .A (sps__n113));
INV_X1 i_0_9_26 (.ZN (n_0_9_25), .A (\mem[1][6] ));
NAND2_X1 i_0_9_25 (.ZN (n_0_9_24), .A1 (n_0_9_34), .A2 (n_0_9_25));
INV_X1 i_0_9_24 (.ZN (n_0_9_23), .A (\mem[9][6] ));
NAND2_X1 i_0_9_23 (.ZN (n_0_9_22), .A1 (sps__n106), .A2 (n_0_9_23));
NAND3_X1 i_0_9_22 (.ZN (n_0_9_21), .A1 (n_0_9_24), .A2 (n_0_9_32), .A3 (n_0_9_22));
NAND3_X1 i_0_9_21 (.ZN (n_0_9_20), .A1 (n_0_9_34), .A2 (\mem[5][6] ), .A3 (address[2]));
NAND3_X1 i_0_9_20 (.ZN (n_0_9_19), .A1 (n_0_9_21), .A2 (n_0_9_26), .A3 (n_0_9_20));
NAND3_X1 i_0_9_19 (.ZN (n_0_9_18), .A1 (n_0_9_19), .A2 (sps__n97), .A3 (n_0_9_27));
INV_X1 i_0_9_18 (.ZN (n_0_9_17), .A (sps__n97));
INV_X1 i_0_9_17 (.ZN (n_0_9_16), .A (\mem[8][6] ));
NAND2_X1 i_0_9_16 (.ZN (n_0_9_15), .A1 (n_0_9_26), .A2 (n_0_9_16));
INV_X1 i_0_9_15 (.ZN (n_0_9_14), .A (\mem[10][6] ));
NAND2_X1 i_0_9_14 (.ZN (n_0_9_13), .A1 (sps__n114), .A2 (n_0_9_14));
NAND3_X1 i_0_9_13 (.ZN (n_0_9_12), .A1 (n_0_9_15), .A2 (n_0_9_32), .A3 (n_0_9_13));
NAND2_X1 i_0_9_12 (.ZN (n_0_9_11), .A1 (n_0_9_12), .A2 (sps__n106));
NAND2_X1 i_0_9_11 (.ZN (n_0_9_10), .A1 (n_0_9_26), .A2 (\mem[0][6] ));
NAND2_X1 i_0_9_10 (.ZN (n_0_9_9), .A1 (sps__n113), .A2 (\mem[2][6] ));
NAND4_X1 i_0_9_9 (.ZN (n_0_9_8), .A1 (n_0_9_10), .A2 (n_0_9_9), .A3 (n_0_9_34), .A4 (n_0_9_32));
NAND2_X1 i_0_9_8 (.ZN (n_0_9_7), .A1 (n_0_9_26), .A2 (\mem[4][6] ));
NAND2_X1 i_0_9_7 (.ZN (n_0_9_6), .A1 (sps__n113), .A2 (\mem[6][6] ));
NAND3_X1 i_0_9_6 (.ZN (n_0_9_5), .A1 (n_0_9_7), .A2 (address[2]), .A3 (n_0_9_6));
NAND4_X1 i_0_9_5 (.ZN (n_0_9_4), .A1 (n_0_9_11), .A2 (n_0_9_17), .A3 (n_0_9_8), .A4 (n_0_9_5));
NAND2_X1 i_0_9_4 (.ZN (n_0_9_3), .A1 (n_0_9_4), .A2 (n_0_9_18));
NAND2_X1 i_0_9_3 (.ZN (n_0_9_2), .A1 (n_0_9_3), .A2 (n_0_5));
INV_X1 i_0_9_2 (.ZN (n_0_9_1), .A (n_0_5));
NAND2_X1 i_0_9_1 (.ZN (n_0_9_0), .A1 (n_0_9_1), .A2 (dataout[6]));
NAND2_X1 i_0_9_0 (.ZN (n_0_15), .A1 (n_0_9_2), .A2 (n_0_9_0));
NAND2_X1 i_0_8_35 (.ZN (n_0_70), .A1 (n_0_8_32), .A2 (n_0_8_34));
NAND2_X1 i_0_8_34 (.ZN (n_0_8_34), .A1 (n_0_8_30), .A2 (n_0_8_33));
NAND2_X1 i_0_8_33 (.ZN (n_0_8_33), .A1 (n_0_8_0), .A2 (n_0_5));
NAND2_X1 i_0_8_31 (.ZN (n_0_8_32), .A1 (n_0_8_30), .A2 (n_0_8_31));
INV_X1 i_0_8_30 (.ZN (n_0_8_31), .A (n_0_8_1));
NAND2_X1 i_0_8_28 (.ZN (n_0_8_30), .A1 (n_0_8_29), .A2 (n_0_8_8));
INV_X1 i_0_8_25 (.ZN (n_0_8_29), .A (n_0_5));
INV_X1 i_0_8_32 (.ZN (n_0_8_8), .A (dataout[8]));
INV_X1 i_0_8_21 (.ZN (n_0_8_28), .A (sps__n99));
NAND2_X1 i_0_8_29 (.ZN (n_0_8_27), .A1 (address[1]), .A2 (\mem[10][8] ));
INV_X1 i_0_8_20 (.ZN (n_0_8_26), .A (address[1]));
NAND2_X1 i_0_8_27 (.ZN (n_0_8_25), .A1 (n_0_8_26), .A2 (\mem[8][8] ));
NAND3_X1 i_0_8_26 (.ZN (n_0_8_24), .A1 (n_0_8_25), .A2 (sps__n104), .A3 (n_0_8_27));
INV_X1 i_0_8_18 (.ZN (n_0_8_23), .A (sps__n104));
NAND2_X1 i_0_8_24 (.ZN (n_0_8_22), .A1 (sps__n112), .A2 (\mem[2][8] ));
NAND2_X1 i_0_8_23 (.ZN (n_0_8_21), .A1 (n_0_8_26), .A2 (\mem[0][8] ));
NAND3_X1 i_0_8_22 (.ZN (n_0_8_20), .A1 (n_0_8_21), .A2 (n_0_8_23), .A3 (n_0_8_22));
NAND2_X1 i_0_8_16 (.ZN (n_0_8_19), .A1 (n_0_8_24), .A2 (n_0_8_20));
NAND2_X1 i_0_8_15 (.ZN (n_0_8_18), .A1 (n_0_8_19), .A2 (n_0_8_28));
INV_X1 i_0_8_19 (.ZN (n_0_8_17), .A (\mem[9][8] ));
NAND2_X1 i_0_8_13 (.ZN (n_0_8_16), .A1 (sps__n104), .A2 (n_0_8_17));
INV_X1 i_0_8_17 (.ZN (n_0_8_15), .A (\mem[1][8] ));
NAND2_X1 i_0_8_12 (.ZN (n_0_8_14), .A1 (n_0_8_23), .A2 (n_0_8_15));
NAND3_X1 i_0_8_11 (.ZN (n_0_8_13), .A1 (n_0_8_14), .A2 (n_0_8_26), .A3 (n_0_8_16));
INV_X1 i_0_8_14 (.ZN (n_0_8_12), .A (\mem[3][8] ));
NOR2_X1 i_0_8_10 (.ZN (n_0_8_11), .A1 (sps__n104), .A2 (n_0_8_12));
AOI21_X1 i_0_8_9 (.ZN (n_0_8_10), .A (n_0_8_28), .B1 (n_0_8_11), .B2 (address[1]));
AOI21_X1 i_0_8_8 (.ZN (n_0_8_9), .A (sps__n122), .B1 (n_0_8_10), .B2 (n_0_8_13));
NAND2_X1 i_0_8_1 (.ZN (n_0_8_1), .A1 (n_0_8_18), .A2 (n_0_8_9));
NAND2_X1 i_0_8_7 (.ZN (n_0_8_7), .A1 (sps__n112), .A2 (\mem[6][8] ));
NAND2_X1 i_0_8_6 (.ZN (n_0_8_6), .A1 (n_0_8_26), .A2 (\mem[4][8] ));
NAND3_X1 i_0_8_5 (.ZN (n_0_8_5), .A1 (n_0_8_6), .A2 (n_0_8_28), .A3 (n_0_8_7));
NAND2_X1 i_0_8_4 (.ZN (n_0_8_4), .A1 (sps__n112), .A2 (\mem[7][8] ));
NAND2_X1 i_0_8_3 (.ZN (n_0_8_3), .A1 (n_0_8_26), .A2 (\mem[5][8] ));
NAND3_X1 i_0_8_2 (.ZN (n_0_8_2), .A1 (n_0_8_3), .A2 (sps__n99), .A3 (n_0_8_4));
NAND4_X1 i_0_8_0 (.ZN (n_0_8_0), .A1 (n_0_8_5), .A2 (n_0_8_2), .A3 (n_0_8_23), .A4 (sps__n122));
INV_X1 i_0_5_37 (.ZN (n_0_5_36), .A (sps__n114));
INV_X1 i_0_5_36 (.ZN (n_0_5_35), .A (sps__n103));
NAND3_X1 i_0_5_35 (.ZN (n_0_5_34), .A1 (n_0_5_35), .A2 (\mem[5][15] ), .A3 (sps__n123));
INV_X1 i_0_5_34 (.ZN (n_0_5_33), .A (sps__n123));
INV_X1 i_0_5_33 (.ZN (n_0_5_32), .A (\mem[1][15] ));
NAND2_X1 i_0_5_32 (.ZN (n_0_5_31), .A1 (n_0_5_35), .A2 (n_0_5_32));
INV_X1 i_0_5_31 (.ZN (n_0_5_30), .A (\mem[9][15] ));
NAND2_X1 i_0_5_30 (.ZN (n_0_5_29), .A1 (sps__n103), .A2 (n_0_5_30));
NAND3_X1 i_0_5_29 (.ZN (n_0_5_28), .A1 (n_0_5_31), .A2 (n_0_5_33), .A3 (n_0_5_29));
NAND3_X1 i_0_5_28 (.ZN (n_0_5_27), .A1 (n_0_5_28), .A2 (n_0_5_36), .A3 (n_0_5_34));
INV_X1 i_0_5_27 (.ZN (n_0_5_26), .A (\mem[3][15] ));
NAND2_X1 i_0_5_26 (.ZN (n_0_5_25), .A1 (n_0_5_33), .A2 (n_0_5_26));
INV_X1 i_0_5_24 (.ZN (n_0_5_24), .A (\mem[7][15] ));
NAND2_X1 i_0_5_23 (.ZN (n_0_5_23), .A1 (sps__n123), .A2 (n_0_5_24));
NAND3_X1 i_0_5_22 (.ZN (n_0_5_22), .A1 (n_0_5_25), .A2 (n_0_5_35), .A3 (n_0_5_23));
NAND2_X1 i_0_5_21 (.ZN (n_0_5_21), .A1 (n_0_5_22), .A2 (sps__n114));
NAND3_X1 i_0_5_20 (.ZN (n_0_5_19), .A1 (n_0_5_27), .A2 (sps__n98), .A3 (n_0_5_21));
INV_X1 i_0_5_19 (.ZN (n_0_5_18), .A (sps__n98));
INV_X1 i_0_5_18 (.ZN (n_0_5_17), .A (\mem[8][15] ));
NAND2_X1 i_0_5_17 (.ZN (n_0_5_16), .A1 (n_0_5_36), .A2 (n_0_5_17));
INV_X1 i_0_5_16 (.ZN (n_0_5_15), .A (\mem[10][15] ));
NAND2_X1 i_0_5_15 (.ZN (n_0_5_14), .A1 (sps__n114), .A2 (n_0_5_15));
NAND3_X1 i_0_5_14 (.ZN (n_0_5_13), .A1 (n_0_5_16), .A2 (n_0_5_33), .A3 (n_0_5_14));
NAND2_X1 i_0_5_13 (.ZN (n_0_5_12), .A1 (n_0_5_13), .A2 (sps__n103));
NAND2_X1 i_0_5_12 (.ZN (n_0_5_11), .A1 (n_0_5_36), .A2 (\mem[0][15] ));
NAND2_X1 i_0_5_11 (.ZN (n_0_5_10), .A1 (sps__n114), .A2 (\mem[2][15] ));
NAND4_X1 i_0_5_10 (.ZN (n_0_5_9), .A1 (n_0_5_11), .A2 (n_0_5_10), .A3 (n_0_5_35), .A4 (n_0_5_33));
NAND2_X1 i_0_5_9 (.ZN (n_0_5_8), .A1 (n_0_5_36), .A2 (\mem[4][15] ));
NAND2_X1 i_0_5_8 (.ZN (n_0_5_7), .A1 (sps__n114), .A2 (\mem[6][15] ));
NAND3_X1 i_0_5_7 (.ZN (n_0_5_6), .A1 (n_0_5_8), .A2 (sps__n123), .A3 (n_0_5_7));
NAND4_X1 i_0_5_6 (.ZN (n_0_5_5), .A1 (n_0_5_12), .A2 (n_0_5_18), .A3 (n_0_5_9), .A4 (n_0_5_6));
NAND2_X1 i_0_5_5 (.ZN (n_0_5_4), .A1 (n_0_5_5), .A2 (n_0_5_19));
NAND2_X1 i_0_5_4 (.ZN (n_0_5_3), .A1 (n_0_5_4), .A2 (n_0_5));
INV_X1 i_0_5_3 (.ZN (n_0_5_2), .A (n_0_5));
INV_X1 i_0_5_2 (.ZN (n_0_5_1), .A (n_0_5_20));
NAND2_X1 i_0_5_1 (.ZN (n_0_5_0), .A1 (n_0_5_2), .A2 (n_0_5_1));
NAND2_X1 i_0_5_0 (.ZN (n_0_69), .A1 (n_0_5_0), .A2 (n_0_5_3));
INV_X1 i_0_5_25 (.ZN (n_0_5_20), .A (dataout[15]));
NAND2_X1 i_0_0_35 (.ZN (n_0_48), .A1 (n_0_0_32), .A2 (n_0_0_34));
NAND2_X1 i_0_0_34 (.ZN (n_0_0_34), .A1 (n_0_0_30), .A2 (n_0_0_33));
NAND2_X1 i_0_0_33 (.ZN (n_0_0_33), .A1 (n_0_0_0), .A2 (n_0_5));
NAND2_X1 i_0_0_31 (.ZN (n_0_0_32), .A1 (n_0_0_30), .A2 (n_0_0_31));
INV_X1 i_0_0_30 (.ZN (n_0_0_31), .A (n_0_0_7));
NAND2_X1 i_0_0_28 (.ZN (n_0_0_30), .A1 (n_0_0_29), .A2 (n_0_0_28));
INV_X1 i_0_0_25 (.ZN (n_0_0_29), .A (n_0_5));
INV_X1 i_0_0_32 (.ZN (n_0_0_28), .A (dataout[7]));
INV_X1 i_0_0_21 (.ZN (n_0_0_27), .A (sps__n99));
NAND2_X1 i_0_0_29 (.ZN (n_0_0_26), .A1 (sps__n112), .A2 (\mem[10][7] ));
INV_X1 i_0_0_20 (.ZN (n_0_0_25), .A (sps__n112));
NAND2_X1 i_0_0_27 (.ZN (n_0_0_24), .A1 (n_0_0_25), .A2 (\mem[8][7] ));
NAND3_X1 i_0_0_26 (.ZN (n_0_0_23), .A1 (n_0_0_24), .A2 (sps__n105), .A3 (n_0_0_26));
INV_X1 i_0_0_18 (.ZN (n_0_0_22), .A (sps__n105));
NAND2_X1 i_0_0_24 (.ZN (n_0_0_21), .A1 (sps__n112), .A2 (\mem[2][7] ));
NAND2_X1 i_0_0_23 (.ZN (n_0_0_20), .A1 (n_0_0_25), .A2 (\mem[0][7] ));
NAND3_X1 i_0_0_22 (.ZN (n_0_0_19), .A1 (n_0_0_20), .A2 (n_0_0_22), .A3 (n_0_0_21));
NAND2_X1 i_0_0_16 (.ZN (n_0_0_18), .A1 (n_0_0_23), .A2 (n_0_0_19));
NAND2_X1 i_0_0_15 (.ZN (n_0_0_17), .A1 (n_0_0_18), .A2 (n_0_0_27));
INV_X1 i_0_0_19 (.ZN (n_0_0_16), .A (\mem[9][7] ));
NAND2_X1 i_0_0_13 (.ZN (n_0_0_15), .A1 (sps__n105), .A2 (n_0_0_16));
INV_X1 i_0_0_17 (.ZN (n_0_0_14), .A (\mem[1][7] ));
NAND2_X1 i_0_0_12 (.ZN (n_0_0_13), .A1 (n_0_0_22), .A2 (n_0_0_14));
NAND3_X1 i_0_0_11 (.ZN (n_0_0_12), .A1 (n_0_0_13), .A2 (n_0_0_25), .A3 (n_0_0_15));
INV_X1 i_0_0_14 (.ZN (n_0_0_11), .A (\mem[3][7] ));
NOR2_X1 i_0_0_10 (.ZN (n_0_0_10), .A1 (sps__n105), .A2 (n_0_0_11));
AOI21_X1 i_0_0_7 (.ZN (n_0_0_9), .A (n_0_0_27), .B1 (n_0_0_10), .B2 (sps__n112));
AOI21_X1 i_0_0_4 (.ZN (n_0_0_8), .A (sps__n122), .B1 (n_0_0_9), .B2 (n_0_0_12));
NAND2_X1 i_0_0_1 (.ZN (n_0_0_7), .A1 (n_0_0_17), .A2 (n_0_0_8));
NAND2_X1 i_0_0_9 (.ZN (n_0_0_6), .A1 (sps__n112), .A2 (\mem[6][7] ));
NAND2_X1 i_0_0_8 (.ZN (n_0_0_5), .A1 (n_0_0_25), .A2 (\mem[4][7] ));
NAND3_X1 i_0_0_3 (.ZN (n_0_0_4), .A1 (n_0_0_5), .A2 (n_0_0_27), .A3 (n_0_0_6));
NAND2_X1 i_0_0_6 (.ZN (n_0_0_3), .A1 (sps__n112), .A2 (\mem[7][7] ));
NAND2_X1 i_0_0_5 (.ZN (n_0_0_2), .A1 (n_0_0_25), .A2 (\mem[5][7] ));
NAND3_X1 i_0_0_2 (.ZN (n_0_0_1), .A1 (n_0_0_2), .A2 (sps__n99), .A3 (n_0_0_3));
NAND4_X1 i_0_0_0 (.ZN (n_0_0_0), .A1 (n_0_0_4), .A2 (n_0_0_1), .A3 (n_0_0_22), .A4 (sps__n122));
DFF_X2 \mem_reg[0][0]  (.Q (\mem[0][0] ), .CK (n_0_32), .D (n_0_7));
DFF_X2 \mem_reg[0][1]  (.Q (\mem[0][1] ), .CK (n_0_32), .D (n_0_184));
DFF_X2 \mem_reg[0][2]  (.Q (\mem[0][2] ), .CK (n_0_32), .D (n_0_179));
DFF_X2 \mem_reg[0][3]  (.Q (\mem[0][3] ), .CK (n_0_32), .D (n_0_178));
DFF_X2 \mem_reg[0][4]  (.Q (\mem[0][4] ), .CK (n_0_32), .D (n_0_177));
DFF_X2 \mem_reg[0][5]  (.Q (\mem[0][5] ), .CK (n_0_32), .D (n_0_157));
DFF_X2 \mem_reg[0][6]  (.Q (\mem[0][6] ), .CK (n_0_32), .D (n_0_144));
DFF_X2 \mem_reg[0][7]  (.Q (\mem[0][7] ), .CK (n_0_32), .D (n_0_133));
DFF_X2 \mem_reg[0][8]  (.Q (\mem[0][8] ), .CK (n_0_32), .D (n_0_122));
DFF_X2 \mem_reg[0][9]  (.Q (\mem[0][9] ), .CK (n_0_32), .D (n_0_109));
DFF_X2 \mem_reg[0][10]  (.Q (\mem[0][10] ), .CK (n_0_32), .D (n_0_96));
DFF_X2 \mem_reg[0][11]  (.Q (\mem[0][11] ), .CK (n_0_32), .D (n_0_85));
DFF_X2 \mem_reg[0][12]  (.Q (\mem[0][12] ), .CK (n_0_32), .D (n_0_64));
DFF_X2 \mem_reg[0][13]  (.Q (\mem[0][13] ), .CK (n_0_32), .D (n_0_53));
DFF_X2 \mem_reg[0][14]  (.Q (\mem[0][14] ), .CK (n_0_32), .D (n_0_40));
DFF_X2 \mem_reg[0][15]  (.Q (\mem[0][15] ), .CK (n_0_32), .D (n_0_27));
DFF_X1 \mem_reg[2][0]  (.Q (\mem[2][0] ), .CK (n_0_32), .D (n_0_196));
DFF_X1 \mem_reg[2][1]  (.Q (\mem[2][1] ), .CK (n_0_32), .D (n_0_182));
DFF_X1 \mem_reg[2][2]  (.Q (\mem[2][2] ), .CK (n_0_32), .D (n_0_173));
DFF_X1 \mem_reg[2][3]  (.Q (\mem[2][3] ), .CK (n_0_32), .D (n_0_172));
DFF_X1 \mem_reg[2][4]  (.Q (\mem[2][4] ), .CK (n_0_32), .D (n_0_171));
DFF_X1 \mem_reg[2][5]  (.Q (\mem[2][5] ), .CK (n_0_32), .D (n_0_155));
DFF_X1 \mem_reg[2][6]  (.Q (\mem[2][6] ), .CK (n_0_32), .D (n_0_142));
DFF_X1 \mem_reg[2][7]  (.Q (\mem[2][7] ), .CK (n_0_32), .D (n_0_131));
DFF_X1 \mem_reg[2][8]  (.Q (\mem[2][8] ), .CK (n_0_32), .D (n_0_120));
DFF_X1 \mem_reg[2][9]  (.Q (\mem[2][9] ), .CK (n_0_32), .D (n_0_107));
DFF_X1 \mem_reg[2][10]  (.Q (\mem[2][10] ), .CK (n_0_32), .D (n_0_94));
DFF_X1 \mem_reg[2][11]  (.Q (\mem[2][11] ), .CK (n_0_32), .D (n_0_83));
DFF_X1 \mem_reg[2][12]  (.Q (\mem[2][12] ), .CK (n_0_32), .D (n_0_62));
DFF_X1 \mem_reg[2][13]  (.Q (\mem[2][13] ), .CK (n_0_32), .D (n_0_51));
DFF_X1 \mem_reg[2][14]  (.Q (\mem[2][14] ), .CK (n_0_32), .D (n_0_38));
DFF_X1 \mem_reg[2][15]  (.Q (\mem[2][15] ), .CK (n_0_32), .D (n_0_25));
DFF_X2 \mem_reg[3][2]  (.Q (\mem[3][2] ), .CK (n_0_32), .D (n_0_3));
DFF_X2 \mem_reg[3][3]  (.Q (\mem[3][3] ), .CK (n_0_32), .D (n_0_193));
DFF_X2 \mem_reg[3][4]  (.Q (\mem[3][4] ), .CK (n_0_32), .D (n_0_170));
DFF_X2 \mem_reg[3][5]  (.Q (\mem[3][5] ), .CK (n_0_32), .D (n_0_154));
DFF_X2 \mem_reg[3][6]  (.Q (\mem[3][6] ), .CK (n_0_32), .D (n_0_141));
DFF_X2 \mem_reg[3][7]  (.Q (\mem[3][7] ), .CK (n_0_32), .D (n_0_130));
DFF_X2 \mem_reg[3][8]  (.Q (\mem[3][8] ), .CK (n_0_32), .D (n_0_119));
DFF_X2 \mem_reg[3][9]  (.Q (\mem[3][9] ), .CK (n_0_32), .D (n_0_106));
DFF_X2 \mem_reg[3][10]  (.Q (\mem[3][10] ), .CK (n_0_32), .D (n_0_93));
DFF_X2 \mem_reg[3][11]  (.Q (\mem[3][11] ), .CK (n_0_32), .D (n_0_82));
DFF_X2 \mem_reg[3][12]  (.Q (\mem[3][12] ), .CK (n_0_32), .D (n_0_61));
DFF_X2 \mem_reg[3][13]  (.Q (\mem[3][13] ), .CK (n_0_32), .D (n_0_50));
DFF_X2 \mem_reg[3][14]  (.Q (\mem[3][14] ), .CK (n_0_32), .D (n_0_37));
DFF_X2 \mem_reg[3][15]  (.Q (\mem[3][15] ), .CK (n_0_32), .D (n_0_24));
INV_X32 i_0_204_0 (.ZN (n_0_32), .A (clk));
INV_X1 i_0_151_2 (.ZN (n_0_151_1), .A (\mem[3][0] ));
NAND2_X1 i_0_151_1 (.ZN (n_0_151_0), .A1 (n_0_116), .A2 (data[0]));
OAI21_X1 i_0_151_0 (.ZN (n_0_14), .A (n_0_151_0), .B1 (n_0_151_1), .B2 (n_0_116));
INV_X1 i_0_117_2 (.ZN (n_0_117_1), .A (\mem[5][0] ));
NAND2_X1 i_0_117_1 (.ZN (n_0_117_0), .A1 (n_0_99), .A2 (data[0]));
OAI21_X1 i_0_117_0 (.ZN (n_0_12), .A (n_0_117_0), .B1 (n_0_117_1), .B2 (n_0_99));
INV_X1 i_0_100_2 (.ZN (n_0_100_1), .A (\mem[6][0] ));
NAND2_X1 i_0_100_1 (.ZN (n_0_100_0), .A1 (n_0_65), .A2 (data[0]));
OAI21_X1 i_0_100_0 (.ZN (n_0_10), .A (n_0_100_0), .B1 (n_0_100_1), .B2 (n_0_65));
NAND2_X1 i_0_192_3 (.ZN (n_0_192_2), .A1 (n_0_67), .A2 (n_0_5));
INV_X1 i_0_192_2 (.ZN (n_0_192_1), .A (n_0_5));
NAND2_X1 i_0_192_1 (.ZN (n_0_192_0), .A1 (n_0_192_1), .A2 (dataout[0]));
NAND2_X1 i_0_192_0 (.ZN (n_0_31), .A1 (n_0_192_2), .A2 (n_0_192_0));
NAND2_X1 i_0_191_3 (.ZN (n_0_191_2), .A1 (n_0_68), .A2 (n_0_5));
INV_X1 i_0_191_2 (.ZN (n_0_191_1), .A (n_0_5));
NAND2_X1 i_0_191_1 (.ZN (n_0_191_0), .A1 (n_0_191_1), .A2 (dataout[1]));
NAND2_X1 i_0_191_0 (.ZN (n_0_13), .A1 (n_0_191_2), .A2 (n_0_191_0));
DFF_X1 \mem_reg[1][0]  (.Q (\mem[1][0] ), .CK (n_0_32), .D (n_0_197));
DFF_X1 \mem_reg[1][1]  (.Q (\mem[1][1] ), .CK (n_0_32), .D (n_0_183));
DFF_X1 \mem_reg[1][2]  (.Q (\mem[1][2] ), .CK (n_0_32), .D (n_0_176));
DFF_X1 \mem_reg[1][3]  (.Q (\mem[1][3] ), .CK (n_0_32), .D (n_0_175));
DFF_X1 \mem_reg[1][4]  (.Q (\mem[1][4] ), .CK (n_0_32), .D (n_0_174));
DFF_X1 \mem_reg[1][5]  (.Q (\mem[1][5] ), .CK (n_0_32), .D (n_0_156));
DFF_X1 \mem_reg[1][6]  (.Q (\mem[1][6] ), .CK (n_0_32), .D (n_0_143));
DFF_X1 \mem_reg[1][7]  (.Q (\mem[1][7] ), .CK (n_0_32), .D (n_0_132));
DFF_X1 \mem_reg[1][8]  (.Q (\mem[1][8] ), .CK (n_0_32), .D (n_0_121));
DFF_X1 \mem_reg[1][9]  (.Q (\mem[1][9] ), .CK (n_0_32), .D (n_0_108));
DFF_X1 \mem_reg[1][10]  (.Q (\mem[1][10] ), .CK (n_0_32), .D (n_0_95));
DFF_X1 \mem_reg[1][11]  (.Q (\mem[1][11] ), .CK (n_0_32), .D (n_0_84));
DFF_X1 \mem_reg[1][12]  (.Q (\mem[1][12] ), .CK (n_0_32), .D (n_0_63));
DFF_X1 \mem_reg[1][13]  (.Q (\mem[1][13] ), .CK (n_0_32), .D (n_0_52));
DFF_X1 \mem_reg[1][14]  (.Q (\mem[1][14] ), .CK (n_0_32), .D (n_0_39));
DFF_X1 \mem_reg[1][15]  (.Q (\mem[1][15] ), .CK (n_0_32), .D (n_0_26));
DFF_X1 \mem_reg[4][0]  (.Q (\mem[4][0] ), .CK (n_0_32), .D (n_0_195));
DFF_X1 \mem_reg[4][1]  (.Q (\mem[4][1] ), .CK (n_0_32), .D (n_0_181));
DFF_X1 \mem_reg[4][2]  (.Q (\mem[4][2] ), .CK (n_0_32), .D (n_0_169));
DFF_X1 \mem_reg[4][3]  (.Q (\mem[4][3] ), .CK (n_0_32), .D (n_0_168));
DFF_X1 \mem_reg[4][4]  (.Q (\mem[4][4] ), .CK (n_0_32), .D (n_0_167));
DFF_X1 \mem_reg[4][5]  (.Q (\mem[4][5] ), .CK (n_0_32), .D (n_0_153));
DFF_X1 \mem_reg[4][6]  (.Q (\mem[4][6] ), .CK (n_0_32), .D (n_0_140));
DFF_X1 \mem_reg[4][7]  (.Q (\mem[4][7] ), .CK (n_0_32), .D (n_0_129));
DFF_X1 \mem_reg[4][8]  (.Q (\mem[4][8] ), .CK (n_0_32), .D (n_0_118));
DFF_X1 \mem_reg[4][9]  (.Q (\mem[4][9] ), .CK (n_0_32), .D (n_0_105));
DFF_X1 \mem_reg[4][10]  (.Q (\mem[4][10] ), .CK (n_0_32), .D (n_0_92));
DFF_X1 \mem_reg[4][11]  (.Q (\mem[4][11] ), .CK (n_0_32), .D (n_0_81));
DFF_X1 \mem_reg[4][12]  (.Q (\mem[4][12] ), .CK (n_0_32), .D (n_0_60));
DFF_X1 \mem_reg[4][13]  (.Q (\mem[4][13] ), .CK (n_0_32), .D (n_0_47));
DFF_X1 \mem_reg[4][14]  (.Q (\mem[4][14] ), .CK (n_0_32), .D (n_0_36));
DFF_X1 \mem_reg[4][15]  (.Q (\mem[4][15] ), .CK (n_0_32), .D (n_0_23));
DFF_X2 \mem_reg[5][2]  (.Q (\mem[5][2] ), .CK (n_0_32), .D (n_0_2));
DFF_X2 \mem_reg[5][3]  (.Q (\mem[5][3] ), .CK (n_0_32), .D (n_0_192));
DFF_X2 \mem_reg[5][4]  (.Q (\mem[5][4] ), .CK (n_0_32), .D (n_0_166));
DFF_X2 \mem_reg[5][5]  (.Q (\mem[5][5] ), .CK (n_0_32), .D (n_0_152));
DFF_X2 \mem_reg[5][6]  (.Q (\mem[5][6] ), .CK (n_0_32), .D (n_0_139));
DFF_X2 \mem_reg[5][7]  (.Q (\mem[5][7] ), .CK (n_0_32), .D (n_0_128));
DFF_X2 \mem_reg[5][8]  (.Q (\mem[5][8] ), .CK (n_0_32), .D (n_0_115));
DFF_X2 \mem_reg[5][9]  (.Q (\mem[5][9] ), .CK (n_0_32), .D (n_0_104));
DFF_X2 \mem_reg[5][10]  (.Q (\mem[5][10] ), .CK (n_0_32), .D (n_0_91));
DFF_X2 \mem_reg[5][11]  (.Q (\mem[5][11] ), .CK (n_0_32), .D (n_0_80));
DFF_X2 \mem_reg[5][12]  (.Q (\mem[5][12] ), .CK (n_0_32), .D (n_0_59));
DFF_X2 \mem_reg[5][13]  (.Q (\mem[5][13] ), .CK (n_0_32), .D (n_0_46));
DFF_X2 \mem_reg[5][14]  (.Q (\mem[5][14] ), .CK (n_0_32), .D (n_0_35));
DFF_X2 \mem_reg[5][15]  (.Q (\mem[5][15] ), .CK (n_0_32), .D (n_0_22));
DFF_X2 \mem_reg[6][2]  (.Q (\mem[6][2] ), .CK (n_0_32), .D (n_0_1));
DFF_X2 \mem_reg[6][3]  (.Q (\mem[6][3] ), .CK (n_0_32), .D (n_0_191));
DFF_X2 \mem_reg[6][4]  (.Q (\mem[6][4] ), .CK (n_0_32), .D (n_0_165));
DFF_X2 \mem_reg[6][5]  (.Q (\mem[6][5] ), .CK (n_0_32), .D (n_0_149));
DFF_X2 \mem_reg[6][6]  (.Q (\mem[6][6] ), .CK (n_0_32), .D (n_0_138));
DFF_X2 \mem_reg[6][7]  (.Q (\mem[6][7] ), .CK (n_0_32), .D (n_0_127));
DFF_X2 \mem_reg[6][8]  (.Q (\mem[6][8] ), .CK (n_0_32), .D (n_0_114));
DFF_X2 \mem_reg[6][9]  (.Q (\mem[6][9] ), .CK (n_0_32), .D (n_0_103));
DFF_X2 \mem_reg[6][10]  (.Q (\mem[6][10] ), .CK (n_0_32), .D (n_0_90));
DFF_X2 \mem_reg[6][11]  (.Q (\mem[6][11] ), .CK (n_0_32), .D (n_0_79));
DFF_X2 \mem_reg[6][12]  (.Q (\mem[6][12] ), .CK (n_0_32), .D (n_0_58));
DFF_X2 \mem_reg[6][13]  (.Q (\mem[6][13] ), .CK (n_0_32), .D (n_0_45));
DFF_X2 \mem_reg[6][14]  (.Q (\mem[6][14] ), .CK (n_0_32), .D (n_0_34));
DFF_X2 \mem_reg[6][15]  (.Q (\mem[6][15] ), .CK (n_0_32), .D (n_0_21));
DFF_X1 \mem_reg[7][0]  (.Q (\mem[7][0] ), .CK (n_0_32), .D (n_0_194));
DFF_X2 \mem_reg[7][1]  (.Q (\mem[7][1] ), .CK (n_0_32), .D (n_0_188));
DFF_X2 \mem_reg[7][2]  (.Q (\mem[7][2] ), .CK (n_0_32), .D (n_0_164));
DFF_X2 \mem_reg[7][3]  (.Q (\mem[7][3] ), .CK (n_0_32), .D (n_0_163));
DFF_X2 \mem_reg[7][4]  (.Q (\mem[7][4] ), .CK (n_0_32), .D (n_0_162));
DFF_X2 \mem_reg[7][5]  (.Q (\mem[7][5] ), .CK (n_0_32), .D (n_0_148));
DFF_X2 \mem_reg[7][6]  (.Q (\mem[7][6] ), .CK (n_0_32), .D (n_0_137));
DFF_X2 \mem_reg[7][7]  (.Q (\mem[7][7] ), .CK (n_0_32), .D (n_0_126));
DFF_X2 \mem_reg[7][8]  (.Q (\mem[7][8] ), .CK (n_0_32), .D (n_0_113));
DFF_X2 \mem_reg[7][9]  (.Q (\mem[7][9] ), .CK (n_0_32), .D (n_0_102));
DFF_X2 \mem_reg[7][10]  (.Q (\mem[7][10] ), .CK (n_0_32), .D (n_0_89));
DFF_X2 \mem_reg[7][11]  (.Q (\mem[7][11] ), .CK (n_0_32), .D (n_0_78));
DFF_X2 \mem_reg[7][12]  (.Q (\mem[7][12] ), .CK (n_0_32), .D (n_0_57));
DFF_X2 \mem_reg[7][13]  (.Q (\mem[7][13] ), .CK (n_0_32), .D (n_0_44));
DFF_X2 \mem_reg[7][14]  (.Q (\mem[7][14] ), .CK (n_0_32), .D (n_0_33));
DFF_X2 \mem_reg[7][15]  (.Q (\mem[7][15] ), .CK (n_0_32), .D (n_0_20));
DFF_X2 \mem_reg[8][0]  (.Q (\mem[8][0] ), .CK (n_0_32), .D (n_0_6));
DFF_X2 \mem_reg[8][1]  (.Q (\mem[8][1] ), .CK (n_0_32), .D (n_0_186));
DFF_X2 \mem_reg[8][2]  (.Q (\mem[8][2] ), .CK (n_0_32), .D (n_0_180));
DFF_X2 \mem_reg[8][3]  (.Q (\mem[8][3] ), .CK (n_0_32), .D (n_0_161));
DFF_X2 \mem_reg[8][4]  (.Q (\mem[8][4] ), .CK (n_0_32), .D (n_0_160));
DFF_X2 \mem_reg[8][5]  (.Q (\mem[8][5] ), .CK (n_0_32), .D (n_0_147));
DFF_X2 \mem_reg[8][6]  (.Q (\mem[8][6] ), .CK (n_0_32), .D (n_0_136));
DFF_X2 \mem_reg[8][7]  (.Q (\mem[8][7] ), .CK (n_0_32), .D (n_0_125));
DFF_X2 \mem_reg[8][8]  (.Q (\mem[8][8] ), .CK (n_0_32), .D (n_0_112));
DFF_X2 \mem_reg[8][9]  (.Q (\mem[8][9] ), .CK (n_0_32), .D (n_0_101));
DFF_X2 \mem_reg[8][10]  (.Q (\mem[8][10] ), .CK (n_0_32), .D (n_0_88));
DFF_X2 \mem_reg[8][11]  (.Q (\mem[8][11] ), .CK (n_0_32), .D (n_0_77));
DFF_X2 \mem_reg[8][12]  (.Q (\mem[8][12] ), .CK (n_0_32), .D (n_0_56));
DFF_X2 \mem_reg[8][13]  (.Q (\mem[8][13] ), .CK (n_0_32), .D (n_0_43));
DFF_X2 \mem_reg[8][14]  (.Q (\mem[8][14] ), .CK (n_0_32), .D (n_0_30));
DFF_X2 \mem_reg[8][15]  (.Q (\mem[8][15] ), .CK (n_0_32), .D (n_0_19));
DFF_X1 \mem_reg[9][0]  (.Q (\mem[9][0] ), .CK (n_0_32), .D (n_0_187));
DFF_X1 \mem_reg[9][1]  (.Q (\mem[9][1] ), .CK (n_0_32), .D (n_0_150));
DFF_X1 \mem_reg[9][2]  (.Q (\mem[9][2] ), .CK (n_0_32), .D (n_0_0));
DFF_X1 \mem_reg[9][3]  (.Q (\mem[9][3] ), .CK (n_0_32), .D (n_0_190));
DFF_X1 \mem_reg[9][4]  (.Q (\mem[9][4] ), .CK (n_0_32), .D (n_0_159));
DFF_X1 \mem_reg[9][5]  (.Q (\mem[9][5] ), .CK (n_0_32), .D (n_0_146));
DFF_X1 \mem_reg[9][6]  (.Q (\mem[9][6] ), .CK (n_0_32), .D (n_0_135));
DFF_X1 \mem_reg[9][7]  (.Q (\mem[9][7] ), .CK (n_0_32), .D (n_0_124));
DFF_X1 \mem_reg[9][8]  (.Q (\mem[9][8] ), .CK (n_0_32), .D (n_0_111));
DFF_X1 \mem_reg[9][9]  (.Q (\mem[9][9] ), .CK (n_0_32), .D (n_0_98));
DFF_X1 \mem_reg[9][10]  (.Q (\mem[9][10] ), .CK (n_0_32), .D (n_0_87));
DFF_X1 \mem_reg[9][11]  (.Q (\mem[9][11] ), .CK (n_0_32), .D (n_0_76));
DFF_X1 \mem_reg[9][12]  (.Q (\mem[9][12] ), .CK (n_0_32), .D (n_0_55));
DFF_X1 \mem_reg[9][13]  (.Q (\mem[9][13] ), .CK (n_0_32), .D (n_0_42));
DFF_X1 \mem_reg[9][14]  (.Q (\mem[9][14] ), .CK (n_0_32), .D (n_0_29));
DFF_X1 \mem_reg[9][15]  (.Q (\mem[9][15] ), .CK (n_0_32), .D (n_0_18));
DFF_X1 \mem_reg[10][0]  (.Q (\mem[10][0] ), .CK (n_0_32), .D (n_0_185));
DFF_X1 \mem_reg[10][1]  (.Q (\mem[10][1] ), .CK (n_0_32), .D (n_0_117));
DFF_X1 \mem_reg[10][2]  (.Q (\mem[10][2] ), .CK (n_0_32), .D (n_0_198));
DFF_X1 \mem_reg[10][3]  (.Q (\mem[10][3] ), .CK (n_0_32), .D (n_0_189));
DFF_X1 \mem_reg[10][4]  (.Q (\mem[10][4] ), .CK (n_0_32), .D (n_0_158));
DFF_X1 \mem_reg[10][5]  (.Q (\mem[10][5] ), .CK (n_0_32), .D (n_0_145));
DFF_X1 \mem_reg[10][6]  (.Q (\mem[10][6] ), .CK (n_0_32), .D (n_0_134));
DFF_X1 \mem_reg[10][7]  (.Q (\mem[10][7] ), .CK (n_0_32), .D (n_0_123));
DFF_X1 \mem_reg[10][8]  (.Q (\mem[10][8] ), .CK (n_0_32), .D (n_0_110));
DFF_X1 \mem_reg[10][9]  (.Q (\mem[10][9] ), .CK (n_0_32), .D (n_0_97));
DFF_X1 \mem_reg[10][10]  (.Q (\mem[10][10] ), .CK (n_0_32), .D (n_0_86));
DFF_X1 \mem_reg[10][11]  (.Q (\mem[10][11] ), .CK (n_0_32), .D (n_0_75));
DFF_X1 \mem_reg[10][12]  (.Q (\mem[10][12] ), .CK (n_0_32), .D (n_0_54));
DFF_X1 \mem_reg[10][13]  (.Q (\mem[10][13] ), .CK (n_0_32), .D (n_0_41));
DFF_X1 \mem_reg[10][14]  (.Q (\mem[10][14] ), .CK (n_0_32), .D (n_0_28));
DFF_X1 \mem_reg[10][15]  (.Q (\mem[10][15] ), .CK (n_0_32), .D (n_0_17));
CLKBUF_X3 sps__L1_c1 (.Z (sps__n1), .A (write_signal));
CLKBUF_X3 sps__L2_c2 (.Z (sps__n2), .A (sps__n1));
CLKBUF_X3 sps__L3_c3 (.Z (sps__n3), .A (sps__n2));
BUF_X4 sps__L1_c7 (.Z (sps__n7), .A (address[13]));
CLKBUF_X3 sps__L2_c8 (.Z (sps__n8), .A (sps__n7));
CLKBUF_X3 sps__L2_c9 (.Z (sps__n9), .A (sps__n7));
CLKBUF_X3 sps__L1_c13 (.Z (sps__n13), .A (address[12]));
CLKBUF_X3 sps__L1_c14 (.Z (sps__n14), .A (address[12]));
CLKBUF_X3 sps__L2_c15 (.Z (sps__n15), .A (sps__n14));
BUF_X4 sps__L1_c19 (.Z (sps__n19), .A (address[5]));
CLKBUF_X3 sps__L1_c20 (.Z (sps__n20), .A (address[5]));
CLKBUF_X3 sps__L2_c21 (.Z (sps__n21), .A (sps__n20));
BUF_X1 sps__L1_c25 (.Z (sps__n25), .A (address[9]));
CLKBUF_X3 sps__L1_c26 (.Z (sps__n26), .A (address[9]));
CLKBUF_X3 sps__L2_c27 (.Z (sps__n27), .A (sps__n26));
BUF_X2 sps__L1_c28 (.Z (sps__n28), .A (address[9]));
INV_X1 sps__L1_c33 (.ZN (sps__n33), .A (address[14]));
INV_X4 sps__L2_c34 (.ZN (sps__n34), .A (sps__n33));
BUF_X1 sps__L3_c35 (.Z (sps__n35), .A (sps__n34));
INV_X4 sps__L2_c36 (.ZN (sps__n36), .A (sps__n33));
BUF_X2 sps__L1_c41 (.Z (sps__n41), .A (address[8]));
CLKBUF_X3 sps__L1_c42 (.Z (sps__n42), .A (address[8]));
BUF_X2 sps__L2_c43 (.Z (sps__n43), .A (sps__n42));
BUF_X2 sps__L2_c44 (.Z (sps__n44), .A (sps__n42));
CLKBUF_X3 sps__L1_c49 (.Z (sps__n49), .A (address[11]));
CLKBUF_X3 sps__L2_c50 (.Z (sps__n50), .A (sps__n49));
CLKBUF_X3 sps__L3_c51 (.Z (sps__n51), .A (sps__n50));
BUF_X4 sps__L1_c55 (.Z (sps__n55), .A (address[10]));
CLKBUF_X3 sps__L2_c56 (.Z (sps__n56), .A (sps__n55));
CLKBUF_X3 sps__L2_c57 (.Z (sps__n57), .A (sps__n55));
CLKBUF_X3 sps__L1_c61 (.Z (sps__n61), .A (RST));
BUF_X4 sps__L2_c62 (.Z (sps__n62), .A (sps__n61));
BUF_X2 sps__L2_c63 (.Z (sps__n63), .A (sps__n61));
CLKBUF_X3 sps__L1_c67 (.Z (sps__n67), .A (address[6]));
CLKBUF_X3 sps__L2_c68 (.Z (sps__n68), .A (sps__n67));
CLKBUF_X3 sps__L3_c69 (.Z (sps__n69), .A (sps__n68));
CLKBUF_X3 sps__L1_c73 (.Z (sps__n73), .A (read_signal));
BUF_X4 sps__L2_c74 (.Z (sps__n74), .A (sps__n73));
CLKBUF_X3 sps__L3_c75 (.Z (sps__n75), .A (sps__n74));
CLKBUF_X3 sps__L1_c79 (.Z (sps__n79), .A (address[4]));
CLKBUF_X3 sps__L1_c80 (.Z (sps__n80), .A (address[4]));
BUF_X4 sps__L2_c81 (.Z (sps__n81), .A (sps__n80));
BUF_X4 sps__L1_c85 (.Z (sps__n85), .A (address[15]));
BUF_X4 sps__L2_c86 (.Z (sps__n86), .A (sps__n85));
CLKBUF_X3 sps__L2_c87 (.Z (sps__n87), .A (sps__n85));
CLKBUF_X3 sps__L1_c91 (.Z (sps__n91), .A (address[7]));
BUF_X4 sps__L1_c92 (.Z (sps__n92), .A (address[7]));
CLKBUF_X3 sps__L1_c93 (.Z (sps__n93), .A (address[7]));
BUF_X4 sps__L1_c97 (.Z (sps__n97), .A (address[0]));
CLKBUF_X3 sps__L2_c98 (.Z (sps__n98), .A (sps__n97));
BUF_X4 sps__L2_c99 (.Z (sps__n99), .A (sps__n97));
BUF_X4 sps__L1_c103 (.Z (sps__n103), .A (address[3]));
BUF_X2 sps__L2_c104 (.Z (sps__n104), .A (sps__n103));
CLKBUF_X3 sps__L2_c105 (.Z (sps__n105), .A (sps__n103));
BUF_X2 sps__L1_c106 (.Z (sps__n106), .A (address[3]));
INV_X1 sps__L1_c111 (.ZN (sps__n111), .A (address[1]));
INV_X8 sps__L2_c112 (.ZN (sps__n112), .A (sps__n111));
BUF_X2 sps__L3_c113 (.Z (sps__n113), .A (sps__n112));
CLKBUF_X3 sps__L4_c114 (.Z (sps__n114), .A (sps__n113));
BUF_X2 sps__L1_c119 (.Z (sps__n119), .A (address[2]));
INV_X1 sps__L1_c120 (.ZN (sps__n120), .A (address[2]));
INV_X4 sps__L2_c121 (.ZN (sps__n121), .A (sps__n120));
CLKBUF_X3 sps__L3_c122 (.Z (sps__n122), .A (sps__n121));
INV_X4 sps__L2_c123 (.ZN (sps__n123), .A (sps__n120));

endmodule //DMA


