module coordinator(clk,RST,interrupt,load,cnn,Din,Dout,ramAddress,ramDataIn,ramDataOut,readSignal,writeSignal);
input clk,RST,interrupt,load,cnn,readSignal,writeSignal;
input[15:0] Din;
output [255:0] Dout;
integer i=0,isLoading=0;
reg[7:0] in1,in2; //should it come from test bench??
input[7:0] ramDataOut,ramDataIn ; //what is ramDataOut
wire [7:0] tempDataToRAM;
reg[31:0] byteIndx;
reg[2:0] bitIndx;
wire[31:0] newByteIndx;
wire[2:0] newBitIndx;
wire doneDecompressHandler;
reg tempWork,tempWorking;
wire ramReadSignal,ramWriteSignal,ramDoneRead,ramDoneWrite,choosedRamWriteSignal;
input[15:0] ramAddress;
reg [7:0] ramDataOutFile,ramDataOutCompressed,ramDataOutToModules;
reg[15:0] ramAdressCompressed,ramAdressFile,ramAdressCnn,tempAdressToRAM;
// test bench => read file image(decompress handler), read 10 files (1-10)
// mux => WriteSignal+1/ReadSignal+1/RamDataIn (coordinator/MUX)
// file handler
// interrupt , stop signal (optional) 

decompress_handler decompress_handler_module(in1,in2,byteIndx,bitIndx,newByteIndx,newBitIndx,tempWork,clk,RST,doneDecompressHandler,tempWorking,ramAdressCompressed,ramDataOutToModules,ramDataOutCompressed,ramReadSignal,ramWriteSignal);
file_handler file_handler_module(load,clk,ramAddress,RST,Din, write,ramAdressFile, ramDataOutFile);
// MUX Write_MUX(ramWriteSignal,selector1);
MUX Data_In_MUX(load,cnn,WriteSignal,ramDataOutCompressed,ramDataOutFile,"00000000",ramDataIn,tempDataToRAM);//make sure of the selectors //done
ST_Bit_MUX Adress_In_MUX(load,cnn,WriteSignal,ramAdressCompressed,ramAdressFile,"00000000",ramAddress,tempAdressToRAM);//make sure of the selectors //done
One_Bit_MUX Write_Mux(load,cnn,WriteSignal,ramWriteSignal,write,"0",writeSignal,choosedRamWriteSignal);// what is 
DMA dma_module(tempAdressToRAM,tempDataToRAM,ramReadSignal,choosedRamWriteSignal,ramDataOutToModules,clk,RST,ramReadSignal,ramWriteSignal);
// MUX Data_Out_MUX(selector0,selector1);
// we may need different ream info for each module that will interact with the ram
always @(clk) begin
   
end

endmodule;