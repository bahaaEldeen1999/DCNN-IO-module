/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed May  5 23:11:33 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2201443790 */

module DMA(address, data, read_signal, write_signal, dataout, clk, RST, doneRead, 
      doneWrite);
   input [15:0]address;
   input [15:0]data;
   input read_signal;
   input write_signal;
   output [15:0]dataout;
   input clk;
   input RST;
   output doneRead;
   output doneWrite;

   wire [15:0]\mem[1] ;
   wire [15:0]\mem[2] ;
   wire [15:0]\mem[3] ;
   wire [15:0]\mem[4] ;
   wire [15:0]\mem[5] ;
   wire [15:0]\mem[6] ;
   wire [15:0]\mem[7] ;
   wire [15:0]\mem[8] ;
   wire [15:0]\mem[9] ;
   wire [15:0]\mem[10] ;
   wire [15:0]\mem[11] ;
   wire [15:0]\mem[12] ;
   wire [15:0]\mem[13] ;
   wire [15:0]\mem[14] ;
   wire [15:0]\mem[15] ;
   wire [15:0]\mem[16] ;
   wire [15:0]\mem[17] ;
   wire [15:0]\mem[18] ;
   wire [15:0]\mem[19] ;
   wire [15:0]\mem[20] ;
   wire [15:0]\mem[21] ;
   wire [15:0]\mem[22] ;
   wire [15:0]\mem[23] ;
   wire [15:0]\mem[24] ;
   wire [15:0]\mem[25] ;
   wire [15:0]\mem[26] ;
   wire [15:0]\mem[27] ;
   wire [15:0]\mem[28] ;
   wire [15:0]\mem[29] ;
   wire [15:0]\mem[30] ;
   wire [15:0]\mem[31] ;
   wire [15:0]\mem[32] ;
   wire [15:0]\mem[33] ;
   wire [15:0]\mem[34] ;
   wire [15:0]\mem[35] ;
   wire [15:0]\mem[36] ;
   wire [15:0]\mem[37] ;
   wire [15:0]\mem[38] ;
   wire [15:0]\mem[39] ;
   wire [15:0]\mem[40] ;
   wire [15:0]\mem[41] ;
   wire [15:0]\mem[42] ;
   wire [15:0]\mem[43] ;
   wire [15:0]\mem[44] ;
   wire [15:0]\mem[45] ;
   wire [15:0]\mem[46] ;
   wire [15:0]\mem[47] ;
   wire [15:0]\mem[48] ;
   wire [15:0]\mem[49] ;
   wire [15:0]\mem[51] ;
   wire [15:0]\mem[50] ;
   wire n_0_815;
   wire n_0_814;
   wire n_0_813;
   wire n_0_812;
   wire n_0_811;
   wire n_0_810;
   wire n_0_809;
   wire n_0_808;
   wire n_0_807;
   wire n_0_806;
   wire n_0_805;
   wire n_0_804;
   wire n_0_803;
   wire n_0_802;
   wire n_0_801;
   wire n_0_800;
   wire n_0_799;
   wire n_0_798;
   wire n_0_797;
   wire n_0_796;
   wire n_0_795;
   wire n_0_794;
   wire n_0_793;
   wire n_0_792;
   wire n_0_791;
   wire n_0_790;
   wire n_0_789;
   wire n_0_788;
   wire n_0_787;
   wire n_0_786;
   wire n_0_785;
   wire n_0_784;
   wire n_0_783;
   wire n_0_782;
   wire n_0_781;
   wire n_0_780;
   wire n_0_779;
   wire n_0_778;
   wire n_0_777;
   wire n_0_776;
   wire n_0_775;
   wire n_0_774;
   wire n_0_773;
   wire n_0_772;
   wire n_0_771;
   wire n_0_770;
   wire n_0_769;
   wire n_0_768;
   wire n_0_767;
   wire n_0_766;
   wire n_0_765;
   wire n_0_764;
   wire n_0_763;
   wire n_0_762;
   wire n_0_761;
   wire n_0_760;
   wire n_0_759;
   wire n_0_758;
   wire n_0_757;
   wire n_0_756;
   wire n_0_755;
   wire n_0_754;
   wire n_0_753;
   wire n_0_752;
   wire n_0_751;
   wire n_0_750;
   wire n_0_749;
   wire n_0_748;
   wire n_0_747;
   wire n_0_746;
   wire n_0_745;
   wire n_0_744;
   wire n_0_743;
   wire n_0_742;
   wire n_0_741;
   wire n_0_740;
   wire n_0_739;
   wire n_0_738;
   wire n_0_737;
   wire n_0_736;
   wire n_0_735;
   wire n_0_734;
   wire n_0_733;
   wire n_0_732;
   wire n_0_731;
   wire n_0_730;
   wire n_0_729;
   wire n_0_728;
   wire n_0_727;
   wire n_0_726;
   wire n_0_725;
   wire n_0_724;
   wire n_0_723;
   wire n_0_722;
   wire n_0_721;
   wire n_0_720;
   wire n_0_719;
   wire n_0_718;
   wire n_0_717;
   wire n_0_716;
   wire n_0_715;
   wire n_0_714;
   wire n_0_713;
   wire n_0_712;
   wire n_0_711;
   wire n_0_710;
   wire n_0_709;
   wire n_0_708;
   wire n_0_707;
   wire n_0_706;
   wire n_0_705;
   wire n_0_704;
   wire n_0_703;
   wire n_0_702;
   wire n_0_701;
   wire n_0_700;
   wire n_0_699;
   wire n_0_698;
   wire n_0_697;
   wire n_0_696;
   wire n_0_695;
   wire n_0_694;
   wire n_0_693;
   wire n_0_692;
   wire n_0_691;
   wire n_0_690;
   wire n_0_689;
   wire n_0_688;
   wire n_0_687;
   wire n_0_686;
   wire n_0_685;
   wire n_0_684;
   wire n_0_683;
   wire n_0_682;
   wire n_0_681;
   wire n_0_680;
   wire n_0_679;
   wire n_0_678;
   wire n_0_677;
   wire n_0_676;
   wire n_0_675;
   wire n_0_674;
   wire n_0_673;
   wire n_0_672;
   wire n_0_671;
   wire n_0_670;
   wire n_0_669;
   wire n_0_668;
   wire n_0_667;
   wire n_0_666;
   wire n_0_665;
   wire n_0_664;
   wire n_0_663;
   wire n_0_662;
   wire n_0_661;
   wire n_0_660;
   wire n_0_659;
   wire n_0_658;
   wire n_0_657;
   wire n_0_656;
   wire n_0_655;
   wire n_0_654;
   wire n_0_653;
   wire n_0_652;
   wire n_0_651;
   wire n_0_650;
   wire n_0_649;
   wire n_0_648;
   wire n_0_647;
   wire n_0_646;
   wire n_0_645;
   wire n_0_644;
   wire n_0_643;
   wire n_0_642;
   wire n_0_641;
   wire n_0_640;
   wire n_0_639;
   wire n_0_638;
   wire n_0_637;
   wire n_0_636;
   wire n_0_635;
   wire n_0_634;
   wire n_0_633;
   wire n_0_632;
   wire n_0_631;
   wire n_0_630;
   wire n_0_629;
   wire n_0_628;
   wire n_0_627;
   wire n_0_626;
   wire n_0_625;
   wire n_0_624;
   wire n_0_623;
   wire n_0_622;
   wire n_0_621;
   wire n_0_620;
   wire n_0_619;
   wire n_0_618;
   wire n_0_617;
   wire n_0_616;
   wire n_0_615;
   wire n_0_614;
   wire n_0_613;
   wire n_0_612;
   wire n_0_611;
   wire n_0_610;
   wire n_0_609;
   wire n_0_608;
   wire n_0_607;
   wire n_0_606;
   wire n_0_605;
   wire n_0_604;
   wire n_0_603;
   wire n_0_602;
   wire n_0_601;
   wire n_0_600;
   wire n_0_599;
   wire n_0_598;
   wire n_0_597;
   wire n_0_596;
   wire n_0_595;
   wire n_0_594;
   wire n_0_593;
   wire n_0_592;
   wire n_0_591;
   wire n_0_590;
   wire n_0_589;
   wire n_0_588;
   wire n_0_587;
   wire n_0_586;
   wire n_0_585;
   wire n_0_584;
   wire n_0_583;
   wire n_0_582;
   wire n_0_581;
   wire n_0_580;
   wire n_0_579;
   wire n_0_578;
   wire n_0_577;
   wire n_0_576;
   wire n_0_575;
   wire n_0_574;
   wire n_0_573;
   wire n_0_572;
   wire n_0_571;
   wire n_0_570;
   wire n_0_569;
   wire n_0_568;
   wire n_0_567;
   wire n_0_566;
   wire n_0_565;
   wire n_0_564;
   wire n_0_563;
   wire n_0_562;
   wire n_0_561;
   wire n_0_560;
   wire n_0_559;
   wire n_0_558;
   wire n_0_557;
   wire n_0_556;
   wire n_0_555;
   wire n_0_554;
   wire n_0_553;
   wire n_0_552;
   wire n_0_551;
   wire n_0_550;
   wire n_0_549;
   wire n_0_548;
   wire n_0_547;
   wire n_0_546;
   wire n_0_545;
   wire n_0_544;
   wire n_0_543;
   wire n_0_542;
   wire n_0_541;
   wire n_0_540;
   wire n_0_539;
   wire n_0_538;
   wire n_0_537;
   wire n_0_536;
   wire n_0_535;
   wire n_0_534;
   wire n_0_533;
   wire n_0_532;
   wire n_0_531;
   wire n_0_530;
   wire n_0_529;
   wire n_0_528;
   wire n_0_527;
   wire n_0_526;
   wire n_0_525;
   wire n_0_524;
   wire n_0_523;
   wire n_0_522;
   wire n_0_521;
   wire n_0_520;
   wire n_0_519;
   wire n_0_518;
   wire n_0_517;
   wire n_0_516;
   wire n_0_515;
   wire n_0_514;
   wire n_0_513;
   wire n_0_512;
   wire n_0_511;
   wire n_0_510;
   wire n_0_509;
   wire n_0_508;
   wire n_0_507;
   wire n_0_506;
   wire n_0_505;
   wire n_0_504;
   wire n_0_503;
   wire n_0_502;
   wire n_0_501;
   wire n_0_500;
   wire n_0_499;
   wire n_0_498;
   wire n_0_497;
   wire n_0_496;
   wire n_0_495;
   wire n_0_494;
   wire n_0_493;
   wire n_0_492;
   wire n_0_491;
   wire n_0_490;
   wire n_0_489;
   wire n_0_488;
   wire n_0_487;
   wire n_0_486;
   wire n_0_485;
   wire n_0_484;
   wire n_0_483;
   wire n_0_482;
   wire n_0_481;
   wire n_0_480;
   wire n_0_479;
   wire n_0_478;
   wire n_0_477;
   wire n_0_476;
   wire n_0_475;
   wire n_0_474;
   wire n_0_473;
   wire n_0_472;
   wire n_0_471;
   wire n_0_470;
   wire n_0_469;
   wire n_0_468;
   wire n_0_467;
   wire n_0_466;
   wire n_0_465;
   wire n_0_464;
   wire n_0_463;
   wire n_0_462;
   wire n_0_461;
   wire n_0_460;
   wire n_0_459;
   wire n_0_458;
   wire n_0_457;
   wire n_0_456;
   wire n_0_455;
   wire n_0_454;
   wire n_0_453;
   wire n_0_452;
   wire n_0_451;
   wire n_0_450;
   wire n_0_449;
   wire n_0_448;
   wire n_0_447;
   wire n_0_446;
   wire n_0_445;
   wire n_0_444;
   wire n_0_443;
   wire n_0_442;
   wire n_0_441;
   wire n_0_440;
   wire n_0_439;
   wire n_0_438;
   wire n_0_437;
   wire n_0_436;
   wire n_0_435;
   wire n_0_434;
   wire n_0_433;
   wire n_0_432;
   wire n_0_431;
   wire n_0_430;
   wire n_0_429;
   wire n_0_428;
   wire n_0_427;
   wire n_0_426;
   wire n_0_425;
   wire n_0_424;
   wire n_0_423;
   wire n_0_422;
   wire n_0_421;
   wire n_0_420;
   wire n_0_419;
   wire n_0_418;
   wire n_0_417;
   wire n_0_416;
   wire n_0_415;
   wire n_0_414;
   wire n_0_413;
   wire n_0_412;
   wire n_0_411;
   wire n_0_410;
   wire n_0_409;
   wire n_0_408;
   wire n_0_407;
   wire n_0_406;
   wire n_0_405;
   wire n_0_404;
   wire n_0_403;
   wire n_0_402;
   wire n_0_401;
   wire n_0_400;
   wire n_0_399;
   wire n_0_398;
   wire n_0_397;
   wire n_0_396;
   wire n_0_395;
   wire n_0_394;
   wire n_0_393;
   wire n_0_392;
   wire n_0_391;
   wire n_0_390;
   wire n_0_389;
   wire n_0_388;
   wire n_0_387;
   wire n_0_386;
   wire n_0_385;
   wire n_0_384;
   wire n_0_383;
   wire n_0_382;
   wire n_0_381;
   wire n_0_380;
   wire n_0_379;
   wire n_0_378;
   wire n_0_377;
   wire n_0_376;
   wire n_0_375;
   wire n_0_374;
   wire n_0_373;
   wire n_0_372;
   wire n_0_371;
   wire n_0_370;
   wire n_0_369;
   wire n_0_368;
   wire n_0_367;
   wire n_0_366;
   wire n_0_365;
   wire n_0_364;
   wire n_0_363;
   wire n_0_362;
   wire n_0_361;
   wire n_0_360;
   wire n_0_359;
   wire n_0_358;
   wire n_0_357;
   wire n_0_356;
   wire n_0_355;
   wire n_0_354;
   wire n_0_353;
   wire n_0_352;
   wire n_0_351;
   wire n_0_350;
   wire n_0_349;
   wire n_0_348;
   wire n_0_347;
   wire n_0_346;
   wire n_0_345;
   wire n_0_344;
   wire n_0_343;
   wire n_0_342;
   wire n_0_341;
   wire n_0_340;
   wire n_0_339;
   wire n_0_338;
   wire n_0_337;
   wire n_0_336;
   wire n_0_335;
   wire n_0_334;
   wire n_0_333;
   wire n_0_332;
   wire n_0_331;
   wire n_0_330;
   wire n_0_329;
   wire n_0_328;
   wire n_0_327;
   wire n_0_326;
   wire n_0_325;
   wire n_0_324;
   wire n_0_323;
   wire n_0_322;
   wire n_0_321;
   wire n_0_320;
   wire n_0_319;
   wire n_0_318;
   wire n_0_317;
   wire n_0_316;
   wire n_0_315;
   wire n_0_314;
   wire n_0_313;
   wire n_0_312;
   wire n_0_311;
   wire n_0_310;
   wire n_0_309;
   wire n_0_308;
   wire n_0_307;
   wire n_0_306;
   wire n_0_305;
   wire n_0_304;
   wire n_0_303;
   wire n_0_302;
   wire n_0_301;
   wire n_0_300;
   wire n_0_299;
   wire n_0_298;
   wire n_0_297;
   wire n_0_296;
   wire n_0_295;
   wire n_0_294;
   wire n_0_293;
   wire n_0_292;
   wire n_0_291;
   wire n_0_290;
   wire n_0_289;
   wire n_0_288;
   wire n_0_287;
   wire n_0_286;
   wire n_0_285;
   wire n_0_284;
   wire n_0_283;
   wire n_0_282;
   wire n_0_281;
   wire n_0_280;
   wire n_0_279;
   wire n_0_278;
   wire n_0_277;
   wire n_0_276;
   wire n_0_275;
   wire n_0_274;
   wire n_0_273;
   wire n_0_272;
   wire n_0_271;
   wire n_0_270;
   wire n_0_269;
   wire n_0_268;
   wire n_0_267;
   wire n_0_266;
   wire n_0_265;
   wire n_0_264;
   wire n_0_263;
   wire n_0_262;
   wire n_0_261;
   wire n_0_260;
   wire n_0_259;
   wire n_0_258;
   wire n_0_257;
   wire n_0_256;
   wire n_0_255;
   wire n_0_254;
   wire n_0_253;
   wire n_0_252;
   wire n_0_251;
   wire n_0_250;
   wire n_0_249;
   wire n_0_248;
   wire n_0_247;
   wire n_0_246;
   wire n_0_245;
   wire n_0_244;
   wire n_0_243;
   wire n_0_242;
   wire n_0_241;
   wire n_0_240;
   wire n_0_239;
   wire n_0_238;
   wire n_0_237;
   wire n_0_236;
   wire n_0_235;
   wire n_0_234;
   wire n_0_233;
   wire n_0_232;
   wire n_0_231;
   wire n_0_230;
   wire n_0_229;
   wire n_0_228;
   wire n_0_227;
   wire n_0_226;
   wire n_0_225;
   wire n_0_224;
   wire n_0_223;
   wire n_0_222;
   wire n_0_221;
   wire n_0_220;
   wire n_0_219;
   wire n_0_218;
   wire n_0_217;
   wire n_0_216;
   wire n_0_215;
   wire n_0_214;
   wire n_0_213;
   wire n_0_212;
   wire n_0_211;
   wire n_0_210;
   wire n_0_209;
   wire n_0_208;
   wire n_0_207;
   wire n_0_206;
   wire n_0_205;
   wire n_0_204;
   wire n_0_203;
   wire n_0_202;
   wire n_0_201;
   wire n_0_200;
   wire n_0_199;
   wire n_0_198;
   wire n_0_197;
   wire n_0_196;
   wire n_0_195;
   wire n_0_194;
   wire n_0_193;
   wire n_0_192;
   wire n_0_191;
   wire n_0_190;
   wire n_0_189;
   wire n_0_188;
   wire n_0_187;
   wire n_0_186;
   wire n_0_185;
   wire n_0_184;
   wire n_0_183;
   wire n_0_182;
   wire n_0_181;
   wire n_0_180;
   wire n_0_179;
   wire n_0_178;
   wire n_0_177;
   wire n_0_176;
   wire n_0_175;
   wire n_0_174;
   wire n_0_173;
   wire n_0_172;
   wire n_0_171;
   wire n_0_170;
   wire n_0_169;
   wire n_0_168;
   wire n_0_167;
   wire n_0_166;
   wire n_0_165;
   wire n_0_164;
   wire n_0_163;
   wire n_0_162;
   wire n_0_161;
   wire n_0_160;
   wire n_0_159;
   wire n_0_158;
   wire n_0_157;
   wire n_0_156;
   wire n_0_155;
   wire n_0_154;
   wire n_0_153;
   wire n_0_152;
   wire n_0_151;
   wire n_0_150;
   wire n_0_149;
   wire n_0_148;
   wire n_0_147;
   wire n_0_146;
   wire n_0_145;
   wire n_0_144;
   wire n_0_143;
   wire n_0_142;
   wire n_0_141;
   wire n_0_140;
   wire n_0_139;
   wire n_0_138;
   wire n_0_137;
   wire n_0_136;
   wire n_0_135;
   wire n_0_134;
   wire n_0_133;
   wire n_0_132;
   wire n_0_131;
   wire n_0_130;
   wire n_0_129;
   wire n_0_128;
   wire n_0_127;
   wire n_0_126;
   wire n_0_125;
   wire n_0_124;
   wire n_0_123;
   wire n_0_122;
   wire n_0_121;
   wire n_0_120;
   wire n_0_119;
   wire n_0_118;
   wire n_0_117;
   wire n_0_116;
   wire n_0_115;
   wire n_0_114;
   wire n_0_113;
   wire n_0_112;
   wire n_0_111;
   wire n_0_110;
   wire n_0_109;
   wire n_0_108;
   wire n_0_107;
   wire n_0_106;
   wire n_0_105;
   wire n_0_104;
   wire n_0_103;
   wire n_0_102;
   wire n_0_101;
   wire n_0_100;
   wire n_0_99;
   wire n_0_98;
   wire n_0_97;
   wire n_0_96;
   wire n_0_95;
   wire n_0_94;
   wire n_0_93;
   wire n_0_92;
   wire n_0_91;
   wire n_0_90;
   wire n_0_89;
   wire n_0_88;
   wire n_0_87;
   wire n_0_86;
   wire n_0_85;
   wire n_0_84;
   wire n_0_83;
   wire n_0_82;
   wire n_0_81;
   wire n_0_80;
   wire n_0_79;
   wire n_0_78;
   wire n_0_77;
   wire n_0_76;
   wire n_0_75;
   wire n_0_74;
   wire n_0_73;
   wire n_0_72;
   wire n_0_71;
   wire n_0_70;
   wire n_0_69;
   wire n_0_68;
   wire n_0_67;
   wire n_0_66;
   wire n_0_65;
   wire n_0_64;
   wire n_0_63;
   wire n_0_62;
   wire n_0_61;
   wire n_0_60;
   wire n_0_59;
   wire n_0_58;
   wire n_0_57;
   wire n_0_56;
   wire n_0_55;
   wire n_0_54;
   wire n_0_53;
   wire n_0_52;
   wire n_0_51;
   wire n_0_50;
   wire n_0_49;
   wire n_0_48;
   wire n_0_47;
   wire n_0_46;
   wire n_0_45;
   wire n_0_44;
   wire n_0_43;
   wire n_0_42;
   wire n_0_41;
   wire n_0_40;
   wire n_0_39;
   wire n_0_38;
   wire n_0_37;
   wire n_0_36;
   wire n_0_35;
   wire n_0_34;
   wire n_0_33;
   wire n_0_32;
   wire n_0_31;
   wire n_0_30;
   wire n_0_29;
   wire n_0_28;
   wire n_0_27;
   wire n_0_26;
   wire n_0_25;
   wire n_0_24;
   wire n_0_23;
   wire n_0_22;
   wire n_0_21;
   wire n_0_20;
   wire n_0_19;
   wire n_0_18;
   wire n_0_17;
   wire n_0_16;
   wire n_0_15;
   wire n_0_14;
   wire n_0_13;
   wire n_0_12;
   wire n_0_11;
   wire n_0_10;
   wire n_0_9;
   wire n_0_8;
   wire n_0_7;
   wire n_0_6;
   wire n_0_5;
   wire n_0_4;
   wire n_0_3;
   wire n_0_2;
   wire n_0_1;
   wire n_0_0;
   wire [15:0]\mem[52] ;
   wire [15:0]\mem[53] ;
   wire [15:0]\mem[54] ;
   wire [15:0]\mem[55] ;
   wire [15:0]\mem[56] ;
   wire [15:0]\mem[57] ;
   wire [15:0]\mem[58] ;
   wire [15:0]\mem[59] ;
   wire [15:0]\mem[60] ;
   wire [15:0]\mem[61] ;
   wire [15:0]\mem[62] ;
   wire [15:0]\mem[63] ;
   wire [15:0]\mem[64] ;
   wire [15:0]\mem[65] ;
   wire [15:0]\mem[66] ;
   wire [15:0]\mem[67] ;
   wire [15:0]\mem[68] ;
   wire [15:0]\mem[69] ;
   wire [15:0]\mem[70] ;
   wire [15:0]\mem[71] ;
   wire [15:0]\mem[72] ;
   wire [15:0]\mem[73] ;
   wire [15:0]\mem[74] ;
   wire [15:0]\mem[75] ;
   wire [15:0]\mem[76] ;
   wire [15:0]\mem[77] ;
   wire [15:0]\mem[78] ;
   wire [15:0]\mem[79] ;
   wire [15:0]\mem[80] ;
   wire [15:0]\mem[81] ;
   wire [15:0]\mem[82] ;
   wire [15:0]\mem[83] ;
   wire [15:0]\mem[84] ;
   wire [15:0]\mem[85] ;
   wire [15:0]\mem[86] ;
   wire [15:0]\mem[87] ;
   wire [15:0]\mem[88] ;
   wire [15:0]\mem[89] ;
   wire [15:0]\mem[90] ;
   wire [15:0]\mem[91] ;
   wire [15:0]\mem[92] ;
   wire [15:0]\mem[93] ;
   wire [15:0]\mem[94] ;
   wire [15:0]\mem[95] ;
   wire [15:0]\mem[96] ;
   wire [15:0]\mem[97] ;
   wire [15:0]\mem[98] ;
   wire [15:0]\mem[99] ;
   wire [15:0]\mem[100] ;
   wire [15:0]\mem[0] ;
   wire n_106_799;
   wire n_106_798;
   wire n_106_797;
   wire n_106_796;
   wire n_106_795;
   wire n_106_794;
   wire n_106_793;
   wire n_106_792;
   wire n_106_791;
   wire n_106_790;
   wire n_106_789;
   wire n_106_788;
   wire n_106_787;
   wire n_106_786;
   wire n_106_785;
   wire n_106_784;
   wire n_106_783;
   wire n_106_782;
   wire n_106_781;
   wire n_106_780;
   wire n_106_779;
   wire n_106_778;
   wire n_106_777;
   wire n_106_776;
   wire n_106_775;
   wire n_106_774;
   wire n_106_773;
   wire n_106_772;
   wire n_106_771;
   wire n_106_770;
   wire n_106_769;
   wire n_106_768;
   wire n_106_767;
   wire n_106_766;
   wire n_106_765;
   wire n_106_764;
   wire n_106_763;
   wire n_106_762;
   wire n_106_761;
   wire n_106_760;
   wire n_106_759;
   wire n_106_758;
   wire n_106_757;
   wire n_106_756;
   wire n_106_755;
   wire n_106_754;
   wire n_106_753;
   wire n_106_752;
   wire n_106_751;
   wire n_106_750;
   wire n_106_749;
   wire n_106_748;
   wire n_106_747;
   wire n_106_746;
   wire n_106_745;
   wire n_106_744;
   wire n_106_743;
   wire n_106_742;
   wire n_106_741;
   wire n_106_740;
   wire n_106_739;
   wire n_106_738;
   wire n_106_737;
   wire n_106_736;
   wire n_106_735;
   wire n_106_734;
   wire n_106_733;
   wire n_106_732;
   wire n_106_731;
   wire n_106_730;
   wire n_106_729;
   wire n_106_728;
   wire n_106_727;
   wire n_106_726;
   wire n_106_725;
   wire n_106_724;
   wire n_106_723;
   wire n_106_722;
   wire n_106_721;
   wire n_106_720;
   wire n_106_719;
   wire n_106_718;
   wire n_106_717;
   wire n_106_716;
   wire n_106_715;
   wire n_106_714;
   wire n_106_713;
   wire n_106_712;
   wire n_106_711;
   wire n_106_710;
   wire n_106_709;
   wire n_106_708;
   wire n_106_707;
   wire n_106_706;
   wire n_106_705;
   wire n_106_704;
   wire n_106_703;
   wire n_106_702;
   wire n_106_701;
   wire n_106_700;
   wire n_106_699;
   wire n_106_698;
   wire n_106_697;
   wire n_106_696;
   wire n_106_695;
   wire n_106_694;
   wire n_106_693;
   wire n_106_692;
   wire n_106_691;
   wire n_106_690;
   wire n_106_689;
   wire n_106_688;
   wire n_106_687;
   wire n_106_686;
   wire n_106_685;
   wire n_106_684;
   wire n_106_683;
   wire n_106_682;
   wire n_106_681;
   wire n_106_680;
   wire n_106_679;
   wire n_106_678;
   wire n_106_677;
   wire n_106_676;
   wire n_106_675;
   wire n_106_674;
   wire n_106_673;
   wire n_106_672;
   wire n_106_671;
   wire n_106_670;
   wire n_106_669;
   wire n_106_668;
   wire n_106_667;
   wire n_106_666;
   wire n_106_665;
   wire n_106_664;
   wire n_106_663;
   wire n_106_662;
   wire n_106_661;
   wire n_106_660;
   wire n_106_659;
   wire n_106_658;
   wire n_106_657;
   wire n_106_656;
   wire n_106_655;
   wire n_106_654;
   wire n_106_653;
   wire n_106_652;
   wire n_106_651;
   wire n_106_650;
   wire n_106_649;
   wire n_106_648;
   wire n_106_647;
   wire n_106_646;
   wire n_106_645;
   wire n_106_644;
   wire n_106_643;
   wire n_106_642;
   wire n_106_641;
   wire n_106_640;
   wire n_106_639;
   wire n_106_638;
   wire n_106_637;
   wire n_106_636;
   wire n_106_635;
   wire n_106_634;
   wire n_106_633;
   wire n_106_632;
   wire n_106_631;
   wire n_106_630;
   wire n_106_629;
   wire n_106_628;
   wire n_106_627;
   wire n_106_626;
   wire n_106_625;
   wire n_106_624;
   wire n_106_623;
   wire n_106_622;
   wire n_106_621;
   wire n_106_620;
   wire n_106_619;
   wire n_106_618;
   wire n_106_617;
   wire n_106_616;
   wire n_106_615;
   wire n_106_614;
   wire n_106_613;
   wire n_106_612;
   wire n_106_611;
   wire n_106_610;
   wire n_106_609;
   wire n_106_608;
   wire n_106_607;
   wire n_106_606;
   wire n_106_605;
   wire n_106_604;
   wire n_106_603;
   wire n_106_602;
   wire n_106_601;
   wire n_106_600;
   wire n_106_599;
   wire n_106_598;
   wire n_106_597;
   wire n_106_596;
   wire n_106_595;
   wire n_106_594;
   wire n_106_593;
   wire n_106_592;
   wire n_106_591;
   wire n_106_590;
   wire n_106_589;
   wire n_106_588;
   wire n_106_587;
   wire n_106_586;
   wire n_106_585;
   wire n_106_584;
   wire n_106_583;
   wire n_106_582;
   wire n_106_581;
   wire n_106_580;
   wire n_106_579;
   wire n_106_578;
   wire n_106_577;
   wire n_106_576;
   wire n_106_575;
   wire n_106_574;
   wire n_106_573;
   wire n_106_572;
   wire n_106_571;
   wire n_106_570;
   wire n_106_569;
   wire n_106_568;
   wire n_106_567;
   wire n_106_566;
   wire n_106_565;
   wire n_106_564;
   wire n_106_563;
   wire n_106_562;
   wire n_106_561;
   wire n_106_560;
   wire n_106_559;
   wire n_106_558;
   wire n_106_557;
   wire n_106_556;
   wire n_106_555;
   wire n_106_554;
   wire n_106_553;
   wire n_106_552;
   wire n_106_551;
   wire n_106_550;
   wire n_106_549;
   wire n_106_548;
   wire n_106_547;
   wire n_106_546;
   wire n_106_545;
   wire n_106_544;
   wire n_106_543;
   wire n_106_542;
   wire n_106_541;
   wire n_106_540;
   wire n_106_539;
   wire n_106_538;
   wire n_106_537;
   wire n_106_536;
   wire n_106_535;
   wire n_106_534;
   wire n_106_533;
   wire n_106_532;
   wire n_106_531;
   wire n_106_530;
   wire n_106_529;
   wire n_106_528;
   wire n_106_527;
   wire n_106_526;
   wire n_106_525;
   wire n_106_524;
   wire n_106_523;
   wire n_106_522;
   wire n_106_521;
   wire n_106_520;
   wire n_106_519;
   wire n_106_518;
   wire n_106_517;
   wire n_106_516;
   wire n_106_515;
   wire n_106_514;
   wire n_106_513;
   wire n_106_512;
   wire n_106_511;
   wire n_106_510;
   wire n_106_509;
   wire n_106_508;
   wire n_106_507;
   wire n_106_506;
   wire n_106_505;
   wire n_106_504;
   wire n_106_503;
   wire n_106_502;
   wire n_106_501;
   wire n_106_500;
   wire n_106_499;
   wire n_106_498;
   wire n_106_497;
   wire n_106_496;
   wire n_106_495;
   wire n_106_494;
   wire n_106_493;
   wire n_106_492;
   wire n_106_491;
   wire n_106_490;
   wire n_106_489;
   wire n_106_488;
   wire n_106_487;
   wire n_106_486;
   wire n_106_485;
   wire n_106_484;
   wire n_106_483;
   wire n_106_482;
   wire n_106_481;
   wire n_106_480;
   wire n_106_479;
   wire n_106_478;
   wire n_106_477;
   wire n_106_476;
   wire n_106_475;
   wire n_106_474;
   wire n_106_473;
   wire n_106_472;
   wire n_106_471;
   wire n_106_470;
   wire n_106_469;
   wire n_106_468;
   wire n_106_467;
   wire n_106_466;
   wire n_106_465;
   wire n_106_464;
   wire n_106_463;
   wire n_106_462;
   wire n_106_461;
   wire n_106_460;
   wire n_106_459;
   wire n_106_458;
   wire n_106_457;
   wire n_106_456;
   wire n_106_455;
   wire n_106_454;
   wire n_106_453;
   wire n_106_452;
   wire n_106_451;
   wire n_106_450;
   wire n_106_449;
   wire n_106_448;
   wire n_106_447;
   wire n_106_446;
   wire n_106_445;
   wire n_106_444;
   wire n_106_443;
   wire n_106_442;
   wire n_106_441;
   wire n_106_440;
   wire n_106_439;
   wire n_106_438;
   wire n_106_437;
   wire n_106_436;
   wire n_106_435;
   wire n_106_434;
   wire n_106_433;
   wire n_106_432;
   wire n_106_431;
   wire n_106_430;
   wire n_106_429;
   wire n_106_428;
   wire n_106_427;
   wire n_106_426;
   wire n_106_425;
   wire n_106_424;
   wire n_106_423;
   wire n_106_422;
   wire n_106_421;
   wire n_106_420;
   wire n_106_419;
   wire n_106_418;
   wire n_106_417;
   wire n_106_416;
   wire n_106_415;
   wire n_106_414;
   wire n_106_413;
   wire n_106_412;
   wire n_106_411;
   wire n_106_410;
   wire n_106_409;
   wire n_106_408;
   wire n_106_407;
   wire n_106_406;
   wire n_106_405;
   wire n_106_404;
   wire n_106_403;
   wire n_106_402;
   wire n_106_401;
   wire n_106_400;
   wire n_106_399;
   wire n_106_398;
   wire n_106_397;
   wire n_106_396;
   wire n_106_395;
   wire n_106_394;
   wire n_106_393;
   wire n_106_392;
   wire n_106_391;
   wire n_106_390;
   wire n_106_389;
   wire n_106_388;
   wire n_106_387;
   wire n_106_386;
   wire n_106_385;
   wire n_106_384;
   wire n_106_383;
   wire n_106_382;
   wire n_106_381;
   wire n_106_380;
   wire n_106_379;
   wire n_106_378;
   wire n_106_377;
   wire n_106_376;
   wire n_106_375;
   wire n_106_374;
   wire n_106_373;
   wire n_106_372;
   wire n_106_371;
   wire n_106_370;
   wire n_106_369;
   wire n_106_368;
   wire n_106_367;
   wire n_106_366;
   wire n_106_365;
   wire n_106_364;
   wire n_106_363;
   wire n_106_362;
   wire n_106_361;
   wire n_106_360;
   wire n_106_359;
   wire n_106_358;
   wire n_106_357;
   wire n_106_356;
   wire n_106_355;
   wire n_106_354;
   wire n_106_353;
   wire n_106_352;
   wire n_106_351;
   wire n_106_350;
   wire n_106_349;
   wire n_106_348;
   wire n_106_347;
   wire n_106_346;
   wire n_106_345;
   wire n_106_344;
   wire n_106_343;
   wire n_106_342;
   wire n_106_341;
   wire n_106_340;
   wire n_106_339;
   wire n_106_338;
   wire n_106_337;
   wire n_106_336;
   wire n_106_335;
   wire n_106_334;
   wire n_106_333;
   wire n_106_332;
   wire n_106_331;
   wire n_106_330;
   wire n_106_329;
   wire n_106_328;
   wire n_106_327;
   wire n_106_326;
   wire n_106_325;
   wire n_106_324;
   wire n_106_323;
   wire n_106_322;
   wire n_106_321;
   wire n_106_320;
   wire n_106_319;
   wire n_106_318;
   wire n_106_317;
   wire n_106_316;
   wire n_106_315;
   wire n_106_314;
   wire n_106_313;
   wire n_106_312;
   wire n_106_311;
   wire n_106_310;
   wire n_106_309;
   wire n_106_308;
   wire n_106_307;
   wire n_106_306;
   wire n_106_305;
   wire n_106_304;
   wire n_106_303;
   wire n_106_302;
   wire n_106_301;
   wire n_106_300;
   wire n_106_299;
   wire n_106_298;
   wire n_106_297;
   wire n_106_296;
   wire n_106_295;
   wire n_106_294;
   wire n_106_293;
   wire n_106_292;
   wire n_106_291;
   wire n_106_290;
   wire n_106_289;
   wire n_106_288;
   wire n_106_287;
   wire n_106_286;
   wire n_106_285;
   wire n_106_284;
   wire n_106_283;
   wire n_106_282;
   wire n_106_281;
   wire n_106_280;
   wire n_106_279;
   wire n_106_278;
   wire n_106_277;
   wire n_106_276;
   wire n_106_275;
   wire n_106_274;
   wire n_106_273;
   wire n_106_272;
   wire n_106_271;
   wire n_106_270;
   wire n_106_269;
   wire n_106_268;
   wire n_106_267;
   wire n_106_266;
   wire n_106_265;
   wire n_106_264;
   wire n_106_263;
   wire n_106_262;
   wire n_106_261;
   wire n_106_260;
   wire n_106_259;
   wire n_106_258;
   wire n_106_257;
   wire n_106_256;
   wire n_106_255;
   wire n_106_254;
   wire n_106_253;
   wire n_106_252;
   wire n_106_251;
   wire n_106_250;
   wire n_106_249;
   wire n_106_248;
   wire n_106_247;
   wire n_106_246;
   wire n_106_245;
   wire n_106_244;
   wire n_106_243;
   wire n_106_242;
   wire n_106_241;
   wire n_106_240;
   wire n_106_239;
   wire n_106_238;
   wire n_106_237;
   wire n_106_236;
   wire n_106_235;
   wire n_106_234;
   wire n_106_233;
   wire n_106_232;
   wire n_106_231;
   wire n_106_230;
   wire n_106_229;
   wire n_106_228;
   wire n_106_227;
   wire n_106_226;
   wire n_106_225;
   wire n_106_224;
   wire n_106_223;
   wire n_106_222;
   wire n_106_221;
   wire n_106_220;
   wire n_106_219;
   wire n_106_218;
   wire n_106_217;
   wire n_106_216;
   wire n_106_215;
   wire n_106_214;
   wire n_106_213;
   wire n_106_212;
   wire n_106_211;
   wire n_106_210;
   wire n_106_209;
   wire n_106_208;
   wire n_106_207;
   wire n_106_206;
   wire n_106_205;
   wire n_106_204;
   wire n_106_203;
   wire n_106_202;
   wire n_106_201;
   wire n_106_200;
   wire n_106_199;
   wire n_106_198;
   wire n_106_197;
   wire n_106_196;
   wire n_106_195;
   wire n_106_194;
   wire n_106_193;
   wire n_106_192;
   wire n_106_191;
   wire n_106_190;
   wire n_106_189;
   wire n_106_188;
   wire n_106_187;
   wire n_106_186;
   wire n_106_185;
   wire n_106_184;
   wire n_106_183;
   wire n_106_182;
   wire n_106_181;
   wire n_106_180;
   wire n_106_179;
   wire n_106_178;
   wire n_106_177;
   wire n_106_176;
   wire n_106_175;
   wire n_106_174;
   wire n_106_173;
   wire n_106_172;
   wire n_106_171;
   wire n_106_170;
   wire n_106_169;
   wire n_106_168;
   wire n_106_167;
   wire n_106_166;
   wire n_106_165;
   wire n_106_164;
   wire n_106_163;
   wire n_106_162;
   wire n_106_161;
   wire n_106_160;
   wire n_106_159;
   wire n_106_158;
   wire n_106_157;
   wire n_106_156;
   wire n_106_155;
   wire n_106_154;
   wire n_106_153;
   wire n_106_152;
   wire n_106_151;
   wire n_106_150;
   wire n_106_149;
   wire n_106_148;
   wire n_106_147;
   wire n_106_146;
   wire n_106_145;
   wire n_106_144;
   wire n_106_143;
   wire n_106_142;
   wire n_106_141;
   wire n_106_140;
   wire n_106_139;
   wire n_106_138;
   wire n_106_137;
   wire n_106_136;
   wire n_106_135;
   wire n_106_134;
   wire n_106_133;
   wire n_106_132;
   wire n_106_131;
   wire n_106_130;
   wire n_106_129;
   wire n_106_128;
   wire n_106_127;
   wire n_106_126;
   wire n_106_125;
   wire n_106_124;
   wire n_106_123;
   wire n_106_122;
   wire n_106_121;
   wire n_106_120;
   wire n_106_119;
   wire n_106_118;
   wire n_106_117;
   wire n_106_116;
   wire n_106_115;
   wire n_106_114;
   wire n_106_113;
   wire n_106_112;
   wire n_106_111;
   wire n_106_110;
   wire n_106_109;
   wire n_106_108;
   wire n_106_107;
   wire n_106_106;
   wire n_106_105;
   wire n_106_104;
   wire n_106_103;
   wire n_106_102;
   wire n_106_101;
   wire n_106_100;
   wire n_106_99;
   wire n_106_98;
   wire n_106_97;
   wire n_106_96;
   wire n_106_95;
   wire n_106_94;
   wire n_106_93;
   wire n_106_92;
   wire n_106_91;
   wire n_106_90;
   wire n_106_89;
   wire n_106_88;
   wire n_106_87;
   wire n_106_86;
   wire n_106_85;
   wire n_106_84;
   wire n_106_83;
   wire n_106_82;
   wire n_106_81;
   wire n_106_80;
   wire n_106_79;
   wire n_106_78;
   wire n_106_77;
   wire n_106_76;
   wire n_106_75;
   wire n_106_74;
   wire n_106_73;
   wire n_106_72;
   wire n_106_71;
   wire n_106_70;
   wire n_106_69;
   wire n_106_68;
   wire n_106_67;
   wire n_106_66;
   wire n_106_65;
   wire n_106_64;
   wire n_106_63;
   wire n_106_62;
   wire n_106_61;
   wire n_106_60;
   wire n_106_59;
   wire n_106_58;
   wire n_106_57;
   wire n_106_56;
   wire n_106_55;
   wire n_106_54;
   wire n_106_53;
   wire n_106_52;
   wire n_106_51;
   wire n_106_50;
   wire n_106_49;
   wire n_106_48;
   wire n_106_47;
   wire n_106_46;
   wire n_106_45;
   wire n_106_44;
   wire n_106_43;
   wire n_106_42;
   wire n_106_41;
   wire n_106_40;
   wire n_106_39;
   wire n_106_38;
   wire n_106_37;
   wire n_106_36;
   wire n_106_35;
   wire n_106_34;
   wire n_106_33;
   wire n_106_32;
   wire n_106_31;
   wire n_106_30;
   wire n_106_29;
   wire n_106_28;
   wire n_106_27;
   wire n_106_26;
   wire n_106_25;
   wire n_106_24;
   wire n_106_23;
   wire n_106_22;
   wire n_106_21;
   wire n_106_20;
   wire n_106_19;
   wire n_106_18;
   wire n_106_17;
   wire n_106_16;
   wire n_106_15;
   wire n_106_14;
   wire n_106_13;
   wire n_106_12;
   wire n_106_11;
   wire n_106_10;
   wire n_106_9;
   wire n_106_8;
   wire n_106_7;
   wire n_106_6;
   wire n_106_5;
   wire n_106_4;
   wire n_106_3;
   wire n_106_2;
   wire n_106_1;
   wire n_106_0;
   wire n_1_0;
   wire n_1_1_0;
   wire n_1_1_1;
   wire n_1_1_2;
   wire n_1_1_3;
   wire n_1_1_4;
   wire n_1_1_5;
   wire n_1_1_6;
   wire n_1_1_7;
   wire n_1_1_8;
   wire n_1_1_9;
   wire n_1_1_10;
   wire n_1_1_11;
   wire n_1_1_12;
   wire n_1_1_13;
   wire n_1_1_14;
   wire n_1_1_15;
   wire n_1_1_16;
   wire n_1_1_17;
   wire n_1_1_18;
   wire n_1_1_19;
   wire n_1_1_20;
   wire n_1_1_21;
   wire n_1_1_22;
   wire n_1_1_23;
   wire n_1_1_24;
   wire n_1_1_25;
   wire n_1_1_26;
   wire n_1_1_27;
   wire n_1_1_28;
   wire n_1_1_29;
   wire n_1_1_30;
   wire n_1_1_31;
   wire n_1_1_32;
   wire n_1_1_33;
   wire n_1_1_34;
   wire n_1_1_35;
   wire n_1_1_36;
   wire n_1_1_37;
   wire n_1_1_38;
   wire n_1_1_39;
   wire n_1_1_40;
   wire n_1_1_41;
   wire n_1_1_42;
   wire n_1_1_43;
   wire n_1_1_44;
   wire n_1_1_45;
   wire n_1_1_46;
   wire n_1_1_47;
   wire n_1_1_48;
   wire n_1_1_49;
   wire n_1_1_50;
   wire n_1_1_51;
   wire n_1_1_52;
   wire n_1_1_53;
   wire n_1_1_54;
   wire n_1_1_55;
   wire n_1_1_56;
   wire n_1_1_57;
   wire n_1_1_58;
   wire n_1_1_59;
   wire n_1_1_60;
   wire n_1_1_61;
   wire n_1_1_62;
   wire n_1_1_63;
   wire n_1_1_64;
   wire n_1_1_65;
   wire n_1_1;
   wire n_1_1_66;
   wire n_1_1_67;
   wire n_1_1_68;
   wire n_1_1_69;
   wire n_1_1_70;
   wire n_1_1_71;
   wire n_1_1_72;
   wire n_1_1_73;
   wire n_1_1_74;
   wire n_1_1_75;
   wire n_1_1_76;
   wire n_1_1_77;
   wire n_1_1_78;
   wire n_1_1_79;
   wire n_1_1_80;
   wire n_1_1_81;
   wire n_1_1_82;
   wire n_1_1_83;
   wire n_1_1_84;
   wire n_1_1_85;
   wire n_1_1_86;
   wire n_1_1_87;
   wire n_1_1_88;
   wire n_1_1_89;
   wire n_1_1_90;
   wire n_1_1_91;
   wire n_1_1_92;
   wire n_1_1_93;
   wire n_1_1_94;
   wire n_1_1_95;
   wire n_1_1_96;
   wire n_1_1_97;
   wire n_1_1_98;
   wire n_1_1_99;
   wire n_1_1_100;
   wire n_1_1_101;
   wire n_1_1_102;
   wire n_1_1_103;
   wire n_1_1_104;
   wire n_1_1_105;
   wire n_1_1_106;
   wire n_1_1_107;
   wire n_1_1_108;
   wire n_1_1_109;
   wire n_1_1_110;
   wire n_1_1_111;
   wire n_1_1_112;
   wire n_1_1_113;
   wire n_1_1_114;
   wire n_1_1_115;
   wire n_1_1_116;
   wire n_1_1_117;
   wire n_1_1_118;
   wire n_1_1_119;
   wire n_1_1_120;
   wire n_1_1_121;
   wire n_1_1_122;
   wire n_1_1_123;
   wire n_1_1_124;
   wire n_1_1_125;
   wire n_1_1_126;
   wire n_1_1_127;
   wire n_1_1_128;
   wire n_1_1_129;
   wire n_1_1_130;
   wire n_1_2;
   wire n_1_1_131;
   wire n_1_1_132;
   wire n_1_1_133;
   wire n_1_1_134;
   wire n_1_1_135;
   wire n_1_1_136;
   wire n_1_1_137;
   wire n_1_1_138;
   wire n_1_1_139;
   wire n_1_1_140;
   wire n_1_1_141;
   wire n_1_1_142;
   wire n_1_1_143;
   wire n_1_1_144;
   wire n_1_1_145;
   wire n_1_1_146;
   wire n_1_1_147;
   wire n_1_1_148;
   wire n_1_1_149;
   wire n_1_1_150;
   wire n_1_1_151;
   wire n_1_1_152;
   wire n_1_1_153;
   wire n_1_1_154;
   wire n_1_1_155;
   wire n_1_1_156;
   wire n_1_1_157;
   wire n_1_1_158;
   wire n_1_1_159;
   wire n_1_1_160;
   wire n_1_1_161;
   wire n_1_1_162;
   wire n_1_1_163;
   wire n_1_1_164;
   wire n_1_1_165;
   wire n_1_1_166;
   wire n_1_1_167;
   wire n_1_1_168;
   wire n_1_1_169;
   wire n_1_1_170;
   wire n_1_1_171;
   wire n_1_1_172;
   wire n_1_1_173;
   wire n_1_1_174;
   wire n_1_1_175;
   wire n_1_1_176;
   wire n_1_1_177;
   wire n_1_1_178;
   wire n_1_1_179;
   wire n_1_1_180;
   wire n_1_1_181;
   wire n_1_1_182;
   wire n_1_1_183;
   wire n_1_1_184;
   wire n_1_1_185;
   wire n_1_1_186;
   wire n_1_1_187;
   wire n_1_1_188;
   wire n_1_1_189;
   wire n_1_1_190;
   wire n_1_1_191;
   wire n_1_1_192;
   wire n_1_3;
   wire n_1_1_193;
   wire n_1_1_194;
   wire n_1_1_195;
   wire n_1_1_196;
   wire n_1_1_197;
   wire n_1_1_198;
   wire n_1_1_199;
   wire n_1_1_200;
   wire n_1_1_201;
   wire n_1_1_202;
   wire n_1_1_203;
   wire n_1_1_204;
   wire n_1_1_205;
   wire n_1_1_206;
   wire n_1_1_207;
   wire n_1_1_208;
   wire n_1_1_209;
   wire n_1_1_210;
   wire n_1_1_211;
   wire n_1_1_212;
   wire n_1_1_213;
   wire n_1_1_214;
   wire n_1_1_215;
   wire n_1_1_216;
   wire n_1_1_217;
   wire n_1_1_218;
   wire n_1_1_219;
   wire n_1_1_220;
   wire n_1_1_221;
   wire n_1_1_222;
   wire n_1_1_223;
   wire n_1_1_224;
   wire n_1_1_225;
   wire n_1_1_226;
   wire n_1_1_227;
   wire n_1_1_228;
   wire n_1_1_229;
   wire n_1_1_230;
   wire n_1_1_231;
   wire n_1_1_232;
   wire n_1_1_233;
   wire n_1_1_234;
   wire n_1_1_235;
   wire n_1_1_236;
   wire n_1_1_237;
   wire n_1_1_238;
   wire n_1_1_239;
   wire n_1_1_240;
   wire n_1_1_241;
   wire n_1_1_242;
   wire n_1_1_243;
   wire n_1_1_244;
   wire n_1_1_245;
   wire n_1_1_246;
   wire n_1_1_247;
   wire n_1_1_248;
   wire n_1_1_249;
   wire n_1_1_250;
   wire n_1_1_251;
   wire n_1_1_252;
   wire n_1_1_253;
   wire n_1_4;
   wire n_1_1_254;
   wire n_1_1_255;
   wire n_1_1_256;
   wire n_1_1_257;
   wire n_1_1_258;
   wire n_1_1_259;
   wire n_1_1_260;
   wire n_1_1_261;
   wire n_1_1_262;
   wire n_1_1_263;
   wire n_1_1_264;
   wire n_1_1_265;
   wire n_1_1_266;
   wire n_1_1_267;
   wire n_1_1_268;
   wire n_1_1_269;
   wire n_1_1_270;
   wire n_1_1_271;
   wire n_1_1_272;
   wire n_1_1_273;
   wire n_1_1_274;
   wire n_1_1_275;
   wire n_1_1_276;
   wire n_1_1_277;
   wire n_1_1_278;
   wire n_1_1_279;
   wire n_1_1_280;
   wire n_1_1_281;
   wire n_1_1_282;
   wire n_1_1_283;
   wire n_1_1_284;
   wire n_1_1_285;
   wire n_1_1_286;
   wire n_1_1_287;
   wire n_1_1_288;
   wire n_1_1_289;
   wire n_1_1_290;
   wire n_1_1_291;
   wire n_1_1_292;
   wire n_1_1_293;
   wire n_1_1_294;
   wire n_1_1_295;
   wire n_1_1_296;
   wire n_1_1_297;
   wire n_1_1_298;
   wire n_1_1_299;
   wire n_1_1_300;
   wire n_1_1_301;
   wire n_1_1_302;
   wire n_1_1_303;
   wire n_1_1_304;
   wire n_1_1_305;
   wire n_1_1_306;
   wire n_1_1_307;
   wire n_1_1_308;
   wire n_1_1_309;
   wire n_1_1_310;
   wire n_1_1_311;
   wire n_1_1_312;
   wire n_1_1_313;
   wire n_1_1_314;
   wire n_1_1_315;
   wire n_1_1_316;
   wire n_1_1_317;
   wire n_1_1_318;
   wire n_1_1_319;
   wire n_1_1_320;
   wire n_1_1_321;
   wire n_1_5;
   wire n_1_1_322;
   wire n_1_1_323;
   wire n_1_1_324;
   wire n_1_1_325;
   wire n_1_1_326;
   wire n_1_1_327;
   wire n_1_1_328;
   wire n_1_1_329;
   wire n_1_1_330;
   wire n_1_1_331;
   wire n_1_1_332;
   wire n_1_1_333;
   wire n_1_1_334;
   wire n_1_1_335;
   wire n_1_1_336;
   wire n_1_1_337;
   wire n_1_1_338;
   wire n_1_1_339;
   wire n_1_1_340;
   wire n_1_1_341;
   wire n_1_1_342;
   wire n_1_1_343;
   wire n_1_1_344;
   wire n_1_1_345;
   wire n_1_1_346;
   wire n_1_1_347;
   wire n_1_1_348;
   wire n_1_1_349;
   wire n_1_1_350;
   wire n_1_1_351;
   wire n_1_1_352;
   wire n_1_1_353;
   wire n_1_1_354;
   wire n_1_1_355;
   wire n_1_1_356;
   wire n_1_1_357;
   wire n_1_1_358;
   wire n_1_1_359;
   wire n_1_1_360;
   wire n_1_1_361;
   wire n_1_1_362;
   wire n_1_1_363;
   wire n_1_1_364;
   wire n_1_1_365;
   wire n_1_1_366;
   wire n_1_1_367;
   wire n_1_1_368;
   wire n_1_1_369;
   wire n_1_1_370;
   wire n_1_1_371;
   wire n_1_1_372;
   wire n_1_1_373;
   wire n_1_1_374;
   wire n_1_1_375;
   wire n_1_1_376;
   wire n_1_1_377;
   wire n_1_1_378;
   wire n_1_1_379;
   wire n_1_1_380;
   wire n_1_1_381;
   wire n_1_1_382;
   wire n_1_1_383;
   wire n_1_1_384;
   wire n_1_6;
   wire n_1_1_385;
   wire n_1_1_386;
   wire n_1_1_387;
   wire n_1_1_388;
   wire n_1_1_389;
   wire n_1_1_390;
   wire n_1_1_391;
   wire n_1_1_392;
   wire n_1_1_393;
   wire n_1_1_394;
   wire n_1_1_395;
   wire n_1_1_396;
   wire n_1_1_397;
   wire n_1_1_398;
   wire n_1_1_399;
   wire n_1_1_400;
   wire n_1_1_401;
   wire n_1_1_402;
   wire n_1_1_403;
   wire n_1_1_404;
   wire n_1_1_405;
   wire n_1_1_406;
   wire n_1_1_407;
   wire n_1_1_408;
   wire n_1_1_409;
   wire n_1_1_410;
   wire n_1_1_411;
   wire n_1_1_412;
   wire n_1_1_413;
   wire n_1_1_414;
   wire n_1_1_415;
   wire n_1_1_416;
   wire n_1_1_417;
   wire n_1_1_418;
   wire n_1_1_419;
   wire n_1_1_420;
   wire n_1_1_421;
   wire n_1_1_422;
   wire n_1_1_423;
   wire n_1_1_424;
   wire n_1_1_425;
   wire n_1_1_426;
   wire n_1_1_427;
   wire n_1_1_428;
   wire n_1_1_429;
   wire n_1_1_430;
   wire n_1_1_431;
   wire n_1_1_432;
   wire n_1_1_433;
   wire n_1_1_434;
   wire n_1_1_435;
   wire n_1_1_436;
   wire n_1_1_437;
   wire n_1_1_438;
   wire n_1_1_439;
   wire n_1_1_440;
   wire n_1_1_441;
   wire n_1_1_442;
   wire n_1_1_443;
   wire n_1_1_444;
   wire n_1_1_445;
   wire n_1_1_446;
   wire n_1_1_447;
   wire n_1_1_448;
   wire n_1_1_449;
   wire n_1_7;
   wire n_1_1_450;
   wire n_1_1_451;
   wire n_1_1_452;
   wire n_1_1_453;
   wire n_1_1_454;
   wire n_1_1_455;
   wire n_1_1_456;
   wire n_1_1_457;
   wire n_1_1_458;
   wire n_1_1_459;
   wire n_1_1_460;
   wire n_1_1_461;
   wire n_1_1_462;
   wire n_1_1_463;
   wire n_1_1_464;
   wire n_1_1_465;
   wire n_1_1_466;
   wire n_1_1_467;
   wire n_1_1_468;
   wire n_1_1_469;
   wire n_1_1_470;
   wire n_1_1_471;
   wire n_1_1_472;
   wire n_1_1_473;
   wire n_1_1_474;
   wire n_1_1_475;
   wire n_1_1_476;
   wire n_1_1_477;
   wire n_1_1_478;
   wire n_1_1_479;
   wire n_1_1_480;
   wire n_1_1_481;
   wire n_1_1_482;
   wire n_1_1_483;
   wire n_1_1_484;
   wire n_1_1_485;
   wire n_1_1_486;
   wire n_1_1_487;
   wire n_1_1_488;
   wire n_1_1_489;
   wire n_1_1_490;
   wire n_1_1_491;
   wire n_1_1_492;
   wire n_1_1_493;
   wire n_1_1_494;
   wire n_1_1_495;
   wire n_1_1_496;
   wire n_1_1_497;
   wire n_1_1_498;
   wire n_1_1_499;
   wire n_1_1_500;
   wire n_1_1_501;
   wire n_1_1_502;
   wire n_1_1_503;
   wire n_1_1_504;
   wire n_1_1_505;
   wire n_1_1_506;
   wire n_1_1_507;
   wire n_1_1_508;
   wire n_1_1_509;
   wire n_1_1_510;
   wire n_1_1_511;
   wire n_1_1_512;
   wire n_1_1_513;
   wire n_1_8;
   wire n_1_1_514;
   wire n_1_1_515;
   wire n_1_1_516;
   wire n_1_1_517;
   wire n_1_1_518;
   wire n_1_1_519;
   wire n_1_1_520;
   wire n_1_1_521;
   wire n_1_1_522;
   wire n_1_1_523;
   wire n_1_1_524;
   wire n_1_1_525;
   wire n_1_1_526;
   wire n_1_1_527;
   wire n_1_1_528;
   wire n_1_1_529;
   wire n_1_1_530;
   wire n_1_1_531;
   wire n_1_1_532;
   wire n_1_1_533;
   wire n_1_1_534;
   wire n_1_1_535;
   wire n_1_1_536;
   wire n_1_1_537;
   wire n_1_1_538;
   wire n_1_1_539;
   wire n_1_1_540;
   wire n_1_1_541;
   wire n_1_1_542;
   wire n_1_1_543;
   wire n_1_1_544;
   wire n_1_1_545;
   wire n_1_1_546;
   wire n_1_1_547;
   wire n_1_1_548;
   wire n_1_1_549;
   wire n_1_1_550;
   wire n_1_1_551;
   wire n_1_1_552;
   wire n_1_1_553;
   wire n_1_1_554;
   wire n_1_1_555;
   wire n_1_1_556;
   wire n_1_1_557;
   wire n_1_1_558;
   wire n_1_1_559;
   wire n_1_1_560;
   wire n_1_1_561;
   wire n_1_1_562;
   wire n_1_1_563;
   wire n_1_1_564;
   wire n_1_1_565;
   wire n_1_1_566;
   wire n_1_1_567;
   wire n_1_1_568;
   wire n_1_1_569;
   wire n_1_1_570;
   wire n_1_1_571;
   wire n_1_1_572;
   wire n_1_1_573;
   wire n_1_1_574;
   wire n_1_1_575;
   wire n_1_1_576;
   wire n_1_9;
   wire n_1_1_577;
   wire n_1_1_578;
   wire n_1_1_579;
   wire n_1_1_580;
   wire n_1_1_581;
   wire n_1_1_582;
   wire n_1_1_583;
   wire n_1_1_584;
   wire n_1_1_585;
   wire n_1_1_586;
   wire n_1_1_587;
   wire n_1_1_588;
   wire n_1_1_589;
   wire n_1_1_590;
   wire n_1_1_591;
   wire n_1_1_592;
   wire n_1_1_593;
   wire n_1_1_594;
   wire n_1_1_595;
   wire n_1_1_596;
   wire n_1_1_597;
   wire n_1_1_598;
   wire n_1_1_599;
   wire n_1_1_600;
   wire n_1_1_601;
   wire n_1_1_602;
   wire n_1_1_603;
   wire n_1_1_604;
   wire n_1_1_605;
   wire n_1_1_606;
   wire n_1_1_607;
   wire n_1_1_608;
   wire n_1_1_609;
   wire n_1_1_610;
   wire n_1_1_611;
   wire n_1_1_612;
   wire n_1_1_613;
   wire n_1_1_614;
   wire n_1_1_615;
   wire n_1_1_616;
   wire n_1_1_617;
   wire n_1_1_618;
   wire n_1_1_619;
   wire n_1_1_620;
   wire n_1_1_621;
   wire n_1_1_622;
   wire n_1_1_623;
   wire n_1_1_624;
   wire n_1_1_625;
   wire n_1_1_626;
   wire n_1_1_627;
   wire n_1_1_628;
   wire n_1_1_629;
   wire n_1_1_630;
   wire n_1_1_631;
   wire n_1_1_632;
   wire n_1_1_633;
   wire n_1_1_634;
   wire n_1_1_635;
   wire n_1_1_636;
   wire n_1_1_637;
   wire n_1_1_638;
   wire n_1_1_639;
   wire n_1_1_640;
   wire n_1_10;
   wire n_1_1_641;
   wire n_1_1_642;
   wire n_1_1_643;
   wire n_1_1_644;
   wire n_1_1_645;
   wire n_1_1_646;
   wire n_1_1_647;
   wire n_1_1_648;
   wire n_1_1_649;
   wire n_1_1_650;
   wire n_1_1_651;
   wire n_1_1_652;
   wire n_1_1_653;
   wire n_1_1_654;
   wire n_1_1_655;
   wire n_1_1_656;
   wire n_1_1_657;
   wire n_1_1_658;
   wire n_1_1_659;
   wire n_1_1_660;
   wire n_1_1_661;
   wire n_1_1_662;
   wire n_1_1_663;
   wire n_1_1_664;
   wire n_1_1_665;
   wire n_1_1_666;
   wire n_1_1_667;
   wire n_1_1_668;
   wire n_1_1_669;
   wire n_1_1_670;
   wire n_1_1_671;
   wire n_1_1_672;
   wire n_1_1_673;
   wire n_1_1_674;
   wire n_1_1_675;
   wire n_1_1_676;
   wire n_1_1_677;
   wire n_1_1_678;
   wire n_1_1_679;
   wire n_1_1_680;
   wire n_1_1_681;
   wire n_1_1_682;
   wire n_1_1_683;
   wire n_1_1_684;
   wire n_1_1_685;
   wire n_1_1_686;
   wire n_1_1_687;
   wire n_1_1_688;
   wire n_1_1_689;
   wire n_1_1_690;
   wire n_1_1_691;
   wire n_1_1_692;
   wire n_1_1_693;
   wire n_1_1_694;
   wire n_1_1_695;
   wire n_1_1_696;
   wire n_1_1_697;
   wire n_1_1_698;
   wire n_1_1_699;
   wire n_1_1_700;
   wire n_1_1_701;
   wire n_1_1_702;
   wire n_1_1_703;
   wire n_1_1_704;
   wire n_1_1_705;
   wire n_1_11;
   wire n_1_1_706;
   wire n_1_1_707;
   wire n_1_1_708;
   wire n_1_1_709;
   wire n_1_1_710;
   wire n_1_1_711;
   wire n_1_1_712;
   wire n_1_1_713;
   wire n_1_1_714;
   wire n_1_1_715;
   wire n_1_1_716;
   wire n_1_1_717;
   wire n_1_1_718;
   wire n_1_1_719;
   wire n_1_1_720;
   wire n_1_1_721;
   wire n_1_1_722;
   wire n_1_1_723;
   wire n_1_1_724;
   wire n_1_1_725;
   wire n_1_1_726;
   wire n_1_1_727;
   wire n_1_1_728;
   wire n_1_1_729;
   wire n_1_1_730;
   wire n_1_1_731;
   wire n_1_1_732;
   wire n_1_1_733;
   wire n_1_1_734;
   wire n_1_1_735;
   wire n_1_1_736;
   wire n_1_1_737;
   wire n_1_1_738;
   wire n_1_1_739;
   wire n_1_1_740;
   wire n_1_1_741;
   wire n_1_1_742;
   wire n_1_1_743;
   wire n_1_1_744;
   wire n_1_1_745;
   wire n_1_1_746;
   wire n_1_1_747;
   wire n_1_1_748;
   wire n_1_1_749;
   wire n_1_1_750;
   wire n_1_1_751;
   wire n_1_1_752;
   wire n_1_1_753;
   wire n_1_1_754;
   wire n_1_1_755;
   wire n_1_1_756;
   wire n_1_1_757;
   wire n_1_1_758;
   wire n_1_1_759;
   wire n_1_1_760;
   wire n_1_1_761;
   wire n_1_1_762;
   wire n_1_1_763;
   wire n_1_1_764;
   wire n_1_1_765;
   wire n_1_1_766;
   wire n_1_1_767;
   wire n_1_1_768;
   wire n_1_1_769;
   wire n_1_1_770;
   wire n_1_12;
   wire n_1_1_771;
   wire n_1_1_772;
   wire n_1_1_773;
   wire n_1_1_774;
   wire n_1_1_775;
   wire n_1_1_776;
   wire n_1_1_777;
   wire n_1_1_778;
   wire n_1_1_779;
   wire n_1_1_780;
   wire n_1_1_781;
   wire n_1_1_782;
   wire n_1_1_783;
   wire n_1_1_784;
   wire n_1_1_785;
   wire n_1_1_786;
   wire n_1_1_787;
   wire n_1_1_788;
   wire n_1_1_789;
   wire n_1_1_790;
   wire n_1_1_791;
   wire n_1_1_792;
   wire n_1_1_793;
   wire n_1_1_794;
   wire n_1_1_795;
   wire n_1_1_796;
   wire n_1_1_797;
   wire n_1_1_798;
   wire n_1_1_799;
   wire n_1_1_800;
   wire n_1_1_801;
   wire n_1_1_802;
   wire n_1_1_803;
   wire n_1_1_804;
   wire n_1_1_805;
   wire n_1_1_806;
   wire n_1_1_807;
   wire n_1_1_808;
   wire n_1_1_809;
   wire n_1_1_810;
   wire n_1_1_811;
   wire n_1_1_812;
   wire n_1_1_813;
   wire n_1_1_814;
   wire n_1_1_815;
   wire n_1_1_816;
   wire n_1_1_817;
   wire n_1_1_818;
   wire n_1_1_819;
   wire n_1_1_820;
   wire n_1_1_821;
   wire n_1_1_822;
   wire n_1_1_823;
   wire n_1_1_824;
   wire n_1_1_825;
   wire n_1_1_826;
   wire n_1_1_827;
   wire n_1_1_828;
   wire n_1_1_829;
   wire n_1_1_830;
   wire n_1_1_831;
   wire n_1_1_832;
   wire n_1_13;
   wire n_1_1_833;
   wire n_1_1_834;
   wire n_1_1_835;
   wire n_1_1_836;
   wire n_1_1_837;
   wire n_1_1_838;
   wire n_1_1_839;
   wire n_1_1_840;
   wire n_1_1_841;
   wire n_1_1_842;
   wire n_1_1_843;
   wire n_1_1_844;
   wire n_1_1_845;
   wire n_1_1_846;
   wire n_1_1_847;
   wire n_1_1_848;
   wire n_1_1_849;
   wire n_1_1_850;
   wire n_1_1_851;
   wire n_1_1_852;
   wire n_1_1_853;
   wire n_1_1_854;
   wire n_1_1_855;
   wire n_1_1_856;
   wire n_1_1_857;
   wire n_1_1_858;
   wire n_1_1_859;
   wire n_1_1_860;
   wire n_1_1_861;
   wire n_1_1_862;
   wire n_1_1_863;
   wire n_1_1_864;
   wire n_1_1_865;
   wire n_1_1_866;
   wire n_1_1_867;
   wire n_1_1_868;
   wire n_1_1_869;
   wire n_1_1_870;
   wire n_1_1_871;
   wire n_1_1_872;
   wire n_1_1_873;
   wire n_1_1_874;
   wire n_1_1_875;
   wire n_1_1_876;
   wire n_1_1_877;
   wire n_1_1_878;
   wire n_1_1_879;
   wire n_1_1_880;
   wire n_1_1_881;
   wire n_1_1_882;
   wire n_1_1_883;
   wire n_1_1_884;
   wire n_1_1_885;
   wire n_1_1_886;
   wire n_1_1_887;
   wire n_1_1_888;
   wire n_1_1_889;
   wire n_1_1_890;
   wire n_1_1_891;
   wire n_1_1_892;
   wire n_1_1_893;
   wire n_1_1_894;
   wire n_1_1_895;
   wire n_1_1_896;
   wire n_1_1_897;
   wire n_1_14;
   wire n_1_1_898;
   wire n_1_1_899;
   wire n_1_1_900;
   wire n_1_1_901;
   wire n_1_1_902;
   wire n_1_1_903;
   wire n_1_1_904;
   wire n_1_1_905;
   wire n_1_1_906;
   wire n_1_1_907;
   wire n_1_1_908;
   wire n_1_1_909;
   wire n_1_1_910;
   wire n_1_1_911;
   wire n_1_1_912;
   wire n_1_1_913;
   wire n_1_1_914;
   wire n_1_1_915;
   wire n_1_1_916;
   wire n_1_1_917;
   wire n_1_1_918;
   wire n_1_1_919;
   wire n_1_1_920;
   wire n_1_1_921;
   wire n_1_1_922;
   wire n_1_1_923;
   wire n_1_1_924;
   wire n_1_1_925;
   wire n_1_1_926;
   wire n_1_1_927;
   wire n_1_1_928;
   wire n_1_1_929;
   wire n_1_1_930;
   wire n_1_1_931;
   wire n_1_1_932;
   wire n_1_1_933;
   wire n_1_1_934;
   wire n_1_1_935;
   wire n_1_1_936;
   wire n_1_1_937;
   wire n_1_1_938;
   wire n_1_1_939;
   wire n_1_1_940;
   wire n_1_1_941;
   wire n_1_1_942;
   wire n_1_1_943;
   wire n_1_1_944;
   wire n_1_1_945;
   wire n_1_1_946;
   wire n_1_1_947;
   wire n_1_1_948;
   wire n_1_1_949;
   wire n_1_1_950;
   wire n_1_1_951;
   wire n_1_1_952;
   wire n_1_1_953;
   wire n_1_1_954;
   wire n_1_1_955;
   wire n_1_1_956;
   wire n_1_1_957;
   wire n_1_1_958;
   wire n_1_1_959;
   wire n_1_1_960;
   wire n_1_1_961;
   wire n_1_1_962;
   wire n_1_1_963;
   wire n_1_15;
   wire n_1_1_964;
   wire n_1_1_965;
   wire n_1_1_966;
   wire n_1_1_967;
   wire n_1_1_968;
   wire n_1_1_969;
   wire n_1_1_970;
   wire n_1_1_971;
   wire n_1_1_972;
   wire n_1_1_973;
   wire n_1_1_974;
   wire n_1_1_975;
   wire n_1_1_976;
   wire n_1_1_977;
   wire n_1_1_978;
   wire n_1_1_979;
   wire n_1_1_980;
   wire n_1_1_981;
   wire n_1_1_982;
   wire n_1_1_983;
   wire n_1_1_984;
   wire n_1_1_985;
   wire n_1_1_986;
   wire n_1_1_987;
   wire n_1_1_988;
   wire n_1_1_989;
   wire n_1_1_990;
   wire n_1_1_991;
   wire n_1_1_992;
   wire n_1_1_993;
   wire n_1_1_994;
   wire n_1_1_995;
   wire n_1_1_996;
   wire n_1_1_997;
   wire n_1_1_998;
   wire n_1_1_999;
   wire n_1_1_1000;
   wire n_1_1_1001;
   wire n_1_1_1002;
   wire n_1_1_1003;
   wire n_1_1_1004;
   wire n_1_1_1005;
   wire n_1_1_1006;
   wire n_1_1_1007;
   wire n_1_1_1008;
   wire n_1_1_1009;
   wire n_1_1_1010;
   wire n_1_1_1011;
   wire n_1_1_1012;
   wire n_1_1_1013;
   wire n_1_1_1014;
   wire n_1_1_1015;
   wire n_1_1_1016;
   wire n_1_1_1017;
   wire n_1_1_1018;
   wire n_1_1_1019;
   wire n_1_1_1020;
   wire n_1_1_1021;
   wire n_1_1_1022;
   wire n_1_1_1023;
   wire n_1_1_1024;
   wire n_1_1_1025;
   wire n_1_1_1026;
   wire n_1_1_1027;
   wire n_1_1_1028;
   wire n_1_1_1029;
   wire n_1_1_1030;
   wire n_1_1_1031;
   wire n_1_1_1032;
   wire n_1_1_1033;
   wire n_1_1_1034;
   wire n_1_1_1035;
   wire n_1_1_1036;
   wire n_1_1_1037;
   wire n_1_1_1038;
   wire n_1_1_1039;
   wire n_1_1_1040;
   wire n_1_1_1041;
   wire n_1_1_1042;
   wire n_1_1_1043;
   wire n_1_1_1044;
   wire n_1_1_1045;
   wire n_1_1_1046;
   wire n_1_1_1047;
   wire n_1_1_1048;
   wire n_1_1_1049;
   wire n_1_1_1050;
   wire n_1_1_1051;
   wire n_1_1_1052;
   wire n_1_1_1053;
   wire n_1_1_1054;
   wire n_1_1_1055;
   wire n_1_1_1056;
   wire n_1_1_1057;
   wire n_1_1_1058;
   wire n_1_1_1059;
   wire n_1_1_1060;
   wire n_1_1_1061;
   wire n_1_1_1062;
   wire n_1_1_1063;
   wire n_1_1_1064;
   wire n_1_1_1065;
   wire n_1_1_1066;
   wire n_1_1_1067;
   wire n_1_1_1068;
   wire n_1_1_1069;
   wire n_1_1_1070;
   wire n_1_1_1071;
   wire n_1_1_1072;
   wire n_1_1_1073;
   wire n_1_1_1074;
   wire n_1_1_1075;
   wire n_1_1_1076;
   wire n_1_1_1077;
   wire n_1_1_1078;
   wire n_1_1_1079;
   wire n_1_1_1080;
   wire n_1_1_1081;
   wire n_1_1_1082;
   wire n_1_1_1083;
   wire n_1_1_1084;
   wire n_1_1_1085;
   wire n_1_1_1086;
   wire n_1_1_1087;
   wire n_1_1_1088;
   wire n_1_1_1089;
   wire n_1_1_1090;
   wire n_1_1_1091;
   wire n_1_1_1092;
   wire n_1_1_1093;
   wire n_1_1_1094;
   wire n_1_1_1095;
   wire n_1_1_1096;
   wire n_1_1_1097;
   wire n_1_1_1098;
   wire n_1_1_1099;
   wire n_1_1_1100;
   wire n_1_1_1101;
   wire n_1_1_1102;
   wire n_1_1_1103;
   wire n_1_1_1104;
   wire n_1_1_1105;
   wire n_1_1_1106;
   wire n_1_1_1107;
   wire n_1_1_1108;
   wire n_1_1_1109;
   wire n_1_1_1110;
   wire n_1_1_1111;
   wire n_1_1_1112;
   wire n_1_1_1113;
   wire n_1_1_1114;
   wire n_1_1_1115;
   wire n_1_1_1116;
   wire n_1_1_1117;
   wire n_1_1_1118;
   wire n_1_1_1119;
   wire n_1_1_1120;
   wire n_1_1_1121;
   wire n_1_1_1122;
   wire n_1_1_1123;
   wire n_1_1_1124;
   wire n_1_1_1125;
   wire n_1_1_1126;
   wire n_1_1_1127;
   wire n_1_1_1128;
   wire n_1_1_1129;
   wire n_1_1_1130;
   wire n_1_1_1131;
   wire n_1_1_1132;
   wire n_1_1_1133;
   wire n_1_1_1134;
   wire n_1_1_1135;
   wire n_1_1_1136;
   wire n_1_1_1137;
   wire n_1_1_1138;
   wire n_1_1_1139;
   wire n_1_1_1140;
   wire n_1_1_1141;
   wire n_1_1_1142;
   wire n_1_1_1143;
   wire n_1_1_1144;
   wire n_1_1_1145;
   wire n_1_1_1146;
   wire n_1_1_1147;
   wire n_1_1_1148;
   wire n_1_1_1149;
   wire n_1_1_1150;
   wire n_1_1_1151;
   wire n_1_1_1152;
   wire n_1_1_1153;
   wire n_1_1_1154;
   wire n_1_1_1155;
   wire n_1_1_1156;
   wire n_1_1_1157;
   wire n_1_1_1158;
   wire n_1_1_1159;
   wire n_1_1_1160;
   wire n_1_1_1161;
   wire n_1_1_1162;
   wire n_1_1_1163;
   wire n_1_1_1164;
   wire n_1_1_1165;
   wire n_1_1_1166;
   wire n_1_1_1167;
   wire n_1_1_1168;
   wire n_1_1_1169;
   wire n_1_1_1170;
   wire n_1_1_1171;
   wire n_1_1_1172;
   wire n_1_1_1173;
   wire n_1_1_1174;
   wire n_1_1_1175;
   wire n_1_1_1176;
   wire n_1_1_1177;
   wire n_1_1_1178;
   wire n_1_1_1179;
   wire n_1_1_1180;
   wire n_1_1_1181;
   wire n_1_1_1182;
   wire n_1_1_1183;
   wire n_1_1_1184;
   wire n_1_1_1185;
   wire n_1_1_1186;
   wire n_1_1_1187;
   wire n_1_1_1188;
   wire n_1_1_1189;
   wire n_1_1_1190;

   assign doneRead = 1'b1;
   assign doneWrite = 1'b1;

   DFF_X1 \mem_reg[1][15]  (.D(n_0_815), .CK(n_0), .Q(\mem[1] [15]), .QN());
   DFF_X1 \mem_reg[1][14]  (.D(n_0_814), .CK(n_0), .Q(\mem[1] [14]), .QN());
   DFF_X1 \mem_reg[1][13]  (.D(n_0_813), .CK(n_0), .Q(\mem[1] [13]), .QN());
   DFF_X1 \mem_reg[1][12]  (.D(n_0_812), .CK(n_0), .Q(\mem[1] [12]), .QN());
   DFF_X1 \mem_reg[1][11]  (.D(n_0_811), .CK(n_0), .Q(\mem[1] [11]), .QN());
   DFF_X1 \mem_reg[1][10]  (.D(n_0_810), .CK(n_0), .Q(\mem[1] [10]), .QN());
   DFF_X1 \mem_reg[1][9]  (.D(n_0_809), .CK(n_0), .Q(\mem[1] [9]), .QN());
   DFF_X1 \mem_reg[1][8]  (.D(n_0_808), .CK(n_0), .Q(\mem[1] [8]), .QN());
   DFF_X1 \mem_reg[1][7]  (.D(n_0_807), .CK(n_0), .Q(\mem[1] [7]), .QN());
   DFF_X1 \mem_reg[1][6]  (.D(n_0_806), .CK(n_0), .Q(\mem[1] [6]), .QN());
   DFF_X1 \mem_reg[1][5]  (.D(n_0_805), .CK(n_0), .Q(\mem[1] [5]), .QN());
   DFF_X1 \mem_reg[1][4]  (.D(n_0_804), .CK(n_0), .Q(\mem[1] [4]), .QN());
   DFF_X1 \mem_reg[1][3]  (.D(n_0_803), .CK(n_0), .Q(\mem[1] [3]), .QN());
   DFF_X1 \mem_reg[1][2]  (.D(n_0_802), .CK(n_0), .Q(\mem[1] [2]), .QN());
   DFF_X1 \mem_reg[1][1]  (.D(n_0_801), .CK(n_0), .Q(\mem[1] [1]), .QN());
   DFF_X1 \mem_reg[1][0]  (.D(n_0_800), .CK(n_0), .Q(\mem[1] [0]), .QN());
   DFF_X1 \mem_reg[2][15]  (.D(n_0_799), .CK(n_0), .Q(\mem[2] [15]), .QN());
   DFF_X1 \mem_reg[2][14]  (.D(n_0_798), .CK(n_0), .Q(\mem[2] [14]), .QN());
   DFF_X1 \mem_reg[2][13]  (.D(n_0_797), .CK(n_0), .Q(\mem[2] [13]), .QN());
   DFF_X1 \mem_reg[2][12]  (.D(n_0_796), .CK(n_0), .Q(\mem[2] [12]), .QN());
   DFF_X1 \mem_reg[2][11]  (.D(n_0_795), .CK(n_0), .Q(\mem[2] [11]), .QN());
   DFF_X1 \mem_reg[2][10]  (.D(n_0_794), .CK(n_0), .Q(\mem[2] [10]), .QN());
   DFF_X1 \mem_reg[2][9]  (.D(n_0_793), .CK(n_0), .Q(\mem[2] [9]), .QN());
   DFF_X1 \mem_reg[2][8]  (.D(n_0_792), .CK(n_0), .Q(\mem[2] [8]), .QN());
   DFF_X1 \mem_reg[2][7]  (.D(n_0_791), .CK(n_0), .Q(\mem[2] [7]), .QN());
   DFF_X1 \mem_reg[2][6]  (.D(n_0_790), .CK(n_0), .Q(\mem[2] [6]), .QN());
   DFF_X1 \mem_reg[2][5]  (.D(n_0_789), .CK(n_0), .Q(\mem[2] [5]), .QN());
   DFF_X1 \mem_reg[2][4]  (.D(n_0_788), .CK(n_0), .Q(\mem[2] [4]), .QN());
   DFF_X1 \mem_reg[2][3]  (.D(n_0_787), .CK(n_0), .Q(\mem[2] [3]), .QN());
   DFF_X1 \mem_reg[2][2]  (.D(n_0_786), .CK(n_0), .Q(\mem[2] [2]), .QN());
   DFF_X1 \mem_reg[2][1]  (.D(n_0_785), .CK(n_0), .Q(\mem[2] [1]), .QN());
   DFF_X1 \mem_reg[2][0]  (.D(n_0_784), .CK(n_0), .Q(\mem[2] [0]), .QN());
   DFF_X1 \mem_reg[3][15]  (.D(n_0_783), .CK(n_0), .Q(\mem[3] [15]), .QN());
   DFF_X1 \mem_reg[3][14]  (.D(n_0_782), .CK(n_0), .Q(\mem[3] [14]), .QN());
   DFF_X1 \mem_reg[3][13]  (.D(n_0_781), .CK(n_0), .Q(\mem[3] [13]), .QN());
   DFF_X1 \mem_reg[3][12]  (.D(n_0_780), .CK(n_0), .Q(\mem[3] [12]), .QN());
   DFF_X1 \mem_reg[3][11]  (.D(n_0_779), .CK(n_0), .Q(\mem[3] [11]), .QN());
   DFF_X1 \mem_reg[3][10]  (.D(n_0_778), .CK(n_0), .Q(\mem[3] [10]), .QN());
   DFF_X1 \mem_reg[3][9]  (.D(n_0_777), .CK(n_0), .Q(\mem[3] [9]), .QN());
   DFF_X1 \mem_reg[3][8]  (.D(n_0_776), .CK(n_0), .Q(\mem[3] [8]), .QN());
   DFF_X1 \mem_reg[3][7]  (.D(n_0_775), .CK(n_0), .Q(\mem[3] [7]), .QN());
   DFF_X1 \mem_reg[3][6]  (.D(n_0_774), .CK(n_0), .Q(\mem[3] [6]), .QN());
   DFF_X1 \mem_reg[3][5]  (.D(n_0_773), .CK(n_0), .Q(\mem[3] [5]), .QN());
   DFF_X1 \mem_reg[3][4]  (.D(n_0_772), .CK(n_0), .Q(\mem[3] [4]), .QN());
   DFF_X1 \mem_reg[3][3]  (.D(n_0_771), .CK(n_0), .Q(\mem[3] [3]), .QN());
   DFF_X1 \mem_reg[3][2]  (.D(n_0_770), .CK(n_0), .Q(\mem[3] [2]), .QN());
   DFF_X1 \mem_reg[3][1]  (.D(n_0_769), .CK(n_0), .Q(\mem[3] [1]), .QN());
   DFF_X1 \mem_reg[3][0]  (.D(n_0_768), .CK(n_0), .Q(\mem[3] [0]), .QN());
   DFF_X1 \mem_reg[4][15]  (.D(n_0_767), .CK(n_0), .Q(\mem[4] [15]), .QN());
   DFF_X1 \mem_reg[4][14]  (.D(n_0_766), .CK(n_0), .Q(\mem[4] [14]), .QN());
   DFF_X1 \mem_reg[4][13]  (.D(n_0_765), .CK(n_0), .Q(\mem[4] [13]), .QN());
   DFF_X1 \mem_reg[4][12]  (.D(n_0_764), .CK(n_0), .Q(\mem[4] [12]), .QN());
   DFF_X1 \mem_reg[4][11]  (.D(n_0_763), .CK(n_0), .Q(\mem[4] [11]), .QN());
   DFF_X1 \mem_reg[4][10]  (.D(n_0_762), .CK(n_0), .Q(\mem[4] [10]), .QN());
   DFF_X1 \mem_reg[4][9]  (.D(n_0_761), .CK(n_0), .Q(\mem[4] [9]), .QN());
   DFF_X1 \mem_reg[4][8]  (.D(n_0_760), .CK(n_0), .Q(\mem[4] [8]), .QN());
   DFF_X1 \mem_reg[4][7]  (.D(n_0_759), .CK(n_0), .Q(\mem[4] [7]), .QN());
   DFF_X1 \mem_reg[4][6]  (.D(n_0_758), .CK(n_0), .Q(\mem[4] [6]), .QN());
   DFF_X1 \mem_reg[4][5]  (.D(n_0_757), .CK(n_0), .Q(\mem[4] [5]), .QN());
   DFF_X1 \mem_reg[4][4]  (.D(n_0_756), .CK(n_0), .Q(\mem[4] [4]), .QN());
   DFF_X1 \mem_reg[4][3]  (.D(n_0_755), .CK(n_0), .Q(\mem[4] [3]), .QN());
   DFF_X1 \mem_reg[4][2]  (.D(n_0_754), .CK(n_0), .Q(\mem[4] [2]), .QN());
   DFF_X1 \mem_reg[4][1]  (.D(n_0_753), .CK(n_0), .Q(\mem[4] [1]), .QN());
   DFF_X1 \mem_reg[4][0]  (.D(n_0_752), .CK(n_0), .Q(\mem[4] [0]), .QN());
   DFF_X1 \mem_reg[5][15]  (.D(n_0_751), .CK(n_0), .Q(\mem[5] [15]), .QN());
   DFF_X1 \mem_reg[5][14]  (.D(n_0_750), .CK(n_0), .Q(\mem[5] [14]), .QN());
   DFF_X1 \mem_reg[5][13]  (.D(n_0_749), .CK(n_0), .Q(\mem[5] [13]), .QN());
   DFF_X1 \mem_reg[5][12]  (.D(n_0_748), .CK(n_0), .Q(\mem[5] [12]), .QN());
   DFF_X1 \mem_reg[5][11]  (.D(n_0_747), .CK(n_0), .Q(\mem[5] [11]), .QN());
   DFF_X1 \mem_reg[5][10]  (.D(n_0_746), .CK(n_0), .Q(\mem[5] [10]), .QN());
   DFF_X1 \mem_reg[5][9]  (.D(n_0_745), .CK(n_0), .Q(\mem[5] [9]), .QN());
   DFF_X1 \mem_reg[5][8]  (.D(n_0_744), .CK(n_0), .Q(\mem[5] [8]), .QN());
   DFF_X1 \mem_reg[5][7]  (.D(n_0_743), .CK(n_0), .Q(\mem[5] [7]), .QN());
   DFF_X1 \mem_reg[5][6]  (.D(n_0_742), .CK(n_0), .Q(\mem[5] [6]), .QN());
   DFF_X1 \mem_reg[5][5]  (.D(n_0_741), .CK(n_0), .Q(\mem[5] [5]), .QN());
   DFF_X1 \mem_reg[5][4]  (.D(n_0_740), .CK(n_0), .Q(\mem[5] [4]), .QN());
   DFF_X1 \mem_reg[5][3]  (.D(n_0_739), .CK(n_0), .Q(\mem[5] [3]), .QN());
   DFF_X1 \mem_reg[5][2]  (.D(n_0_738), .CK(n_0), .Q(\mem[5] [2]), .QN());
   DFF_X1 \mem_reg[5][1]  (.D(n_0_737), .CK(n_0), .Q(\mem[5] [1]), .QN());
   DFF_X1 \mem_reg[5][0]  (.D(n_0_736), .CK(n_0), .Q(\mem[5] [0]), .QN());
   DFF_X1 \mem_reg[6][15]  (.D(n_0_735), .CK(n_0), .Q(\mem[6] [15]), .QN());
   DFF_X1 \mem_reg[6][14]  (.D(n_0_734), .CK(n_0), .Q(\mem[6] [14]), .QN());
   DFF_X1 \mem_reg[6][13]  (.D(n_0_733), .CK(n_0), .Q(\mem[6] [13]), .QN());
   DFF_X1 \mem_reg[6][12]  (.D(n_0_732), .CK(n_0), .Q(\mem[6] [12]), .QN());
   DFF_X1 \mem_reg[6][11]  (.D(n_0_731), .CK(n_0), .Q(\mem[6] [11]), .QN());
   DFF_X1 \mem_reg[6][10]  (.D(n_0_730), .CK(n_0), .Q(\mem[6] [10]), .QN());
   DFF_X1 \mem_reg[6][9]  (.D(n_0_729), .CK(n_0), .Q(\mem[6] [9]), .QN());
   DFF_X1 \mem_reg[6][8]  (.D(n_0_728), .CK(n_0), .Q(\mem[6] [8]), .QN());
   DFF_X1 \mem_reg[6][7]  (.D(n_0_727), .CK(n_0), .Q(\mem[6] [7]), .QN());
   DFF_X1 \mem_reg[6][6]  (.D(n_0_726), .CK(n_0), .Q(\mem[6] [6]), .QN());
   DFF_X1 \mem_reg[6][5]  (.D(n_0_725), .CK(n_0), .Q(\mem[6] [5]), .QN());
   DFF_X1 \mem_reg[6][4]  (.D(n_0_724), .CK(n_0), .Q(\mem[6] [4]), .QN());
   DFF_X1 \mem_reg[6][3]  (.D(n_0_723), .CK(n_0), .Q(\mem[6] [3]), .QN());
   DFF_X1 \mem_reg[6][2]  (.D(n_0_722), .CK(n_0), .Q(\mem[6] [2]), .QN());
   DFF_X1 \mem_reg[6][1]  (.D(n_0_721), .CK(n_0), .Q(\mem[6] [1]), .QN());
   DFF_X1 \mem_reg[6][0]  (.D(n_0_720), .CK(n_0), .Q(\mem[6] [0]), .QN());
   DFF_X1 \mem_reg[7][15]  (.D(n_0_719), .CK(n_0), .Q(\mem[7] [15]), .QN());
   DFF_X1 \mem_reg[7][14]  (.D(n_0_718), .CK(n_0), .Q(\mem[7] [14]), .QN());
   DFF_X1 \mem_reg[7][13]  (.D(n_0_717), .CK(n_0), .Q(\mem[7] [13]), .QN());
   DFF_X1 \mem_reg[7][12]  (.D(n_0_716), .CK(n_0), .Q(\mem[7] [12]), .QN());
   DFF_X1 \mem_reg[7][11]  (.D(n_0_715), .CK(n_0), .Q(\mem[7] [11]), .QN());
   DFF_X1 \mem_reg[7][10]  (.D(n_0_714), .CK(n_0), .Q(\mem[7] [10]), .QN());
   DFF_X1 \mem_reg[7][9]  (.D(n_0_713), .CK(n_0), .Q(\mem[7] [9]), .QN());
   DFF_X1 \mem_reg[7][8]  (.D(n_0_712), .CK(n_0), .Q(\mem[7] [8]), .QN());
   DFF_X1 \mem_reg[7][7]  (.D(n_0_711), .CK(n_0), .Q(\mem[7] [7]), .QN());
   DFF_X1 \mem_reg[7][6]  (.D(n_0_710), .CK(n_0), .Q(\mem[7] [6]), .QN());
   DFF_X1 \mem_reg[7][5]  (.D(n_0_709), .CK(n_0), .Q(\mem[7] [5]), .QN());
   DFF_X1 \mem_reg[7][4]  (.D(n_0_708), .CK(n_0), .Q(\mem[7] [4]), .QN());
   DFF_X1 \mem_reg[7][3]  (.D(n_0_707), .CK(n_0), .Q(\mem[7] [3]), .QN());
   DFF_X1 \mem_reg[7][2]  (.D(n_0_706), .CK(n_0), .Q(\mem[7] [2]), .QN());
   DFF_X1 \mem_reg[7][1]  (.D(n_0_705), .CK(n_0), .Q(\mem[7] [1]), .QN());
   DFF_X1 \mem_reg[7][0]  (.D(n_0_704), .CK(n_0), .Q(\mem[7] [0]), .QN());
   DFF_X1 \mem_reg[8][15]  (.D(n_0_703), .CK(n_0), .Q(\mem[8] [15]), .QN());
   DFF_X1 \mem_reg[8][14]  (.D(n_0_702), .CK(n_0), .Q(\mem[8] [14]), .QN());
   DFF_X1 \mem_reg[8][13]  (.D(n_0_701), .CK(n_0), .Q(\mem[8] [13]), .QN());
   DFF_X1 \mem_reg[8][12]  (.D(n_0_700), .CK(n_0), .Q(\mem[8] [12]), .QN());
   DFF_X1 \mem_reg[8][11]  (.D(n_0_699), .CK(n_0), .Q(\mem[8] [11]), .QN());
   DFF_X1 \mem_reg[8][10]  (.D(n_0_698), .CK(n_0), .Q(\mem[8] [10]), .QN());
   DFF_X1 \mem_reg[8][9]  (.D(n_0_697), .CK(n_0), .Q(\mem[8] [9]), .QN());
   DFF_X1 \mem_reg[8][8]  (.D(n_0_696), .CK(n_0), .Q(\mem[8] [8]), .QN());
   DFF_X1 \mem_reg[8][7]  (.D(n_0_695), .CK(n_0), .Q(\mem[8] [7]), .QN());
   DFF_X1 \mem_reg[8][6]  (.D(n_0_694), .CK(n_0), .Q(\mem[8] [6]), .QN());
   DFF_X1 \mem_reg[8][5]  (.D(n_0_693), .CK(n_0), .Q(\mem[8] [5]), .QN());
   DFF_X1 \mem_reg[8][4]  (.D(n_0_692), .CK(n_0), .Q(\mem[8] [4]), .QN());
   DFF_X1 \mem_reg[8][3]  (.D(n_0_691), .CK(n_0), .Q(\mem[8] [3]), .QN());
   DFF_X1 \mem_reg[8][2]  (.D(n_0_690), .CK(n_0), .Q(\mem[8] [2]), .QN());
   DFF_X1 \mem_reg[8][1]  (.D(n_0_689), .CK(n_0), .Q(\mem[8] [1]), .QN());
   DFF_X1 \mem_reg[8][0]  (.D(n_0_688), .CK(n_0), .Q(\mem[8] [0]), .QN());
   DFF_X1 \mem_reg[9][15]  (.D(n_0_687), .CK(n_0), .Q(\mem[9] [15]), .QN());
   DFF_X1 \mem_reg[9][14]  (.D(n_0_686), .CK(n_0), .Q(\mem[9] [14]), .QN());
   DFF_X1 \mem_reg[9][13]  (.D(n_0_685), .CK(n_0), .Q(\mem[9] [13]), .QN());
   DFF_X1 \mem_reg[9][12]  (.D(n_0_684), .CK(n_0), .Q(\mem[9] [12]), .QN());
   DFF_X1 \mem_reg[9][11]  (.D(n_0_683), .CK(n_0), .Q(\mem[9] [11]), .QN());
   DFF_X1 \mem_reg[9][10]  (.D(n_0_682), .CK(n_0), .Q(\mem[9] [10]), .QN());
   DFF_X1 \mem_reg[9][9]  (.D(n_0_681), .CK(n_0), .Q(\mem[9] [9]), .QN());
   DFF_X1 \mem_reg[9][8]  (.D(n_0_680), .CK(n_0), .Q(\mem[9] [8]), .QN());
   DFF_X1 \mem_reg[9][7]  (.D(n_0_679), .CK(n_0), .Q(\mem[9] [7]), .QN());
   DFF_X1 \mem_reg[9][6]  (.D(n_0_678), .CK(n_0), .Q(\mem[9] [6]), .QN());
   DFF_X1 \mem_reg[9][5]  (.D(n_0_677), .CK(n_0), .Q(\mem[9] [5]), .QN());
   DFF_X1 \mem_reg[9][4]  (.D(n_0_676), .CK(n_0), .Q(\mem[9] [4]), .QN());
   DFF_X1 \mem_reg[9][3]  (.D(n_0_675), .CK(n_0), .Q(\mem[9] [3]), .QN());
   DFF_X1 \mem_reg[9][2]  (.D(n_0_674), .CK(n_0), .Q(\mem[9] [2]), .QN());
   DFF_X1 \mem_reg[9][1]  (.D(n_0_673), .CK(n_0), .Q(\mem[9] [1]), .QN());
   DFF_X1 \mem_reg[9][0]  (.D(n_0_672), .CK(n_0), .Q(\mem[9] [0]), .QN());
   DFF_X1 \mem_reg[10][15]  (.D(n_0_671), .CK(n_0), .Q(\mem[10] [15]), .QN());
   DFF_X1 \mem_reg[10][14]  (.D(n_0_670), .CK(n_0), .Q(\mem[10] [14]), .QN());
   DFF_X1 \mem_reg[10][13]  (.D(n_0_669), .CK(n_0), .Q(\mem[10] [13]), .QN());
   DFF_X1 \mem_reg[10][12]  (.D(n_0_668), .CK(n_0), .Q(\mem[10] [12]), .QN());
   DFF_X1 \mem_reg[10][11]  (.D(n_0_667), .CK(n_0), .Q(\mem[10] [11]), .QN());
   DFF_X1 \mem_reg[10][10]  (.D(n_0_666), .CK(n_0), .Q(\mem[10] [10]), .QN());
   DFF_X1 \mem_reg[10][9]  (.D(n_0_665), .CK(n_0), .Q(\mem[10] [9]), .QN());
   DFF_X1 \mem_reg[10][8]  (.D(n_0_664), .CK(n_0), .Q(\mem[10] [8]), .QN());
   DFF_X1 \mem_reg[10][7]  (.D(n_0_663), .CK(n_0), .Q(\mem[10] [7]), .QN());
   DFF_X1 \mem_reg[10][6]  (.D(n_0_662), .CK(n_0), .Q(\mem[10] [6]), .QN());
   DFF_X1 \mem_reg[10][5]  (.D(n_0_661), .CK(n_0), .Q(\mem[10] [5]), .QN());
   DFF_X1 \mem_reg[10][4]  (.D(n_0_660), .CK(n_0), .Q(\mem[10] [4]), .QN());
   DFF_X1 \mem_reg[10][3]  (.D(n_0_659), .CK(n_0), .Q(\mem[10] [3]), .QN());
   DFF_X1 \mem_reg[10][2]  (.D(n_0_658), .CK(n_0), .Q(\mem[10] [2]), .QN());
   DFF_X1 \mem_reg[10][1]  (.D(n_0_657), .CK(n_0), .Q(\mem[10] [1]), .QN());
   DFF_X1 \mem_reg[10][0]  (.D(n_0_656), .CK(n_0), .Q(\mem[10] [0]), .QN());
   DFF_X1 \mem_reg[11][15]  (.D(n_0_655), .CK(n_0), .Q(\mem[11] [15]), .QN());
   DFF_X1 \mem_reg[11][14]  (.D(n_0_654), .CK(n_0), .Q(\mem[11] [14]), .QN());
   DFF_X1 \mem_reg[11][13]  (.D(n_0_653), .CK(n_0), .Q(\mem[11] [13]), .QN());
   DFF_X1 \mem_reg[11][12]  (.D(n_0_652), .CK(n_0), .Q(\mem[11] [12]), .QN());
   DFF_X1 \mem_reg[11][11]  (.D(n_0_651), .CK(n_0), .Q(\mem[11] [11]), .QN());
   DFF_X1 \mem_reg[11][10]  (.D(n_0_650), .CK(n_0), .Q(\mem[11] [10]), .QN());
   DFF_X1 \mem_reg[11][9]  (.D(n_0_649), .CK(n_0), .Q(\mem[11] [9]), .QN());
   DFF_X1 \mem_reg[11][8]  (.D(n_0_648), .CK(n_0), .Q(\mem[11] [8]), .QN());
   DFF_X1 \mem_reg[11][7]  (.D(n_0_647), .CK(n_0), .Q(\mem[11] [7]), .QN());
   DFF_X1 \mem_reg[11][6]  (.D(n_0_646), .CK(n_0), .Q(\mem[11] [6]), .QN());
   DFF_X1 \mem_reg[11][5]  (.D(n_0_645), .CK(n_0), .Q(\mem[11] [5]), .QN());
   DFF_X1 \mem_reg[11][4]  (.D(n_0_644), .CK(n_0), .Q(\mem[11] [4]), .QN());
   DFF_X1 \mem_reg[11][3]  (.D(n_0_643), .CK(n_0), .Q(\mem[11] [3]), .QN());
   DFF_X1 \mem_reg[11][2]  (.D(n_0_642), .CK(n_0), .Q(\mem[11] [2]), .QN());
   DFF_X1 \mem_reg[11][1]  (.D(n_0_641), .CK(n_0), .Q(\mem[11] [1]), .QN());
   DFF_X1 \mem_reg[11][0]  (.D(n_0_640), .CK(n_0), .Q(\mem[11] [0]), .QN());
   DFF_X1 \mem_reg[12][15]  (.D(n_0_639), .CK(n_0), .Q(\mem[12] [15]), .QN());
   DFF_X1 \mem_reg[12][14]  (.D(n_0_638), .CK(n_0), .Q(\mem[12] [14]), .QN());
   DFF_X1 \mem_reg[12][13]  (.D(n_0_637), .CK(n_0), .Q(\mem[12] [13]), .QN());
   DFF_X1 \mem_reg[12][12]  (.D(n_0_636), .CK(n_0), .Q(\mem[12] [12]), .QN());
   DFF_X1 \mem_reg[12][11]  (.D(n_0_635), .CK(n_0), .Q(\mem[12] [11]), .QN());
   DFF_X1 \mem_reg[12][10]  (.D(n_0_634), .CK(n_0), .Q(\mem[12] [10]), .QN());
   DFF_X1 \mem_reg[12][9]  (.D(n_0_633), .CK(n_0), .Q(\mem[12] [9]), .QN());
   DFF_X1 \mem_reg[12][8]  (.D(n_0_632), .CK(n_0), .Q(\mem[12] [8]), .QN());
   DFF_X1 \mem_reg[12][7]  (.D(n_0_631), .CK(n_0), .Q(\mem[12] [7]), .QN());
   DFF_X1 \mem_reg[12][6]  (.D(n_0_630), .CK(n_0), .Q(\mem[12] [6]), .QN());
   DFF_X1 \mem_reg[12][5]  (.D(n_0_629), .CK(n_0), .Q(\mem[12] [5]), .QN());
   DFF_X1 \mem_reg[12][4]  (.D(n_0_628), .CK(n_0), .Q(\mem[12] [4]), .QN());
   DFF_X1 \mem_reg[12][3]  (.D(n_0_627), .CK(n_0), .Q(\mem[12] [3]), .QN());
   DFF_X1 \mem_reg[12][2]  (.D(n_0_626), .CK(n_0), .Q(\mem[12] [2]), .QN());
   DFF_X1 \mem_reg[12][1]  (.D(n_0_625), .CK(n_0), .Q(\mem[12] [1]), .QN());
   DFF_X1 \mem_reg[12][0]  (.D(n_0_624), .CK(n_0), .Q(\mem[12] [0]), .QN());
   DFF_X1 \mem_reg[13][15]  (.D(n_0_623), .CK(n_0), .Q(\mem[13] [15]), .QN());
   DFF_X1 \mem_reg[13][14]  (.D(n_0_622), .CK(n_0), .Q(\mem[13] [14]), .QN());
   DFF_X1 \mem_reg[13][13]  (.D(n_0_621), .CK(n_0), .Q(\mem[13] [13]), .QN());
   DFF_X1 \mem_reg[13][12]  (.D(n_0_620), .CK(n_0), .Q(\mem[13] [12]), .QN());
   DFF_X1 \mem_reg[13][11]  (.D(n_0_619), .CK(n_0), .Q(\mem[13] [11]), .QN());
   DFF_X1 \mem_reg[13][10]  (.D(n_0_618), .CK(n_0), .Q(\mem[13] [10]), .QN());
   DFF_X1 \mem_reg[13][9]  (.D(n_0_617), .CK(n_0), .Q(\mem[13] [9]), .QN());
   DFF_X1 \mem_reg[13][8]  (.D(n_0_616), .CK(n_0), .Q(\mem[13] [8]), .QN());
   DFF_X1 \mem_reg[13][7]  (.D(n_0_615), .CK(n_0), .Q(\mem[13] [7]), .QN());
   DFF_X1 \mem_reg[13][6]  (.D(n_0_614), .CK(n_0), .Q(\mem[13] [6]), .QN());
   DFF_X1 \mem_reg[13][5]  (.D(n_0_613), .CK(n_0), .Q(\mem[13] [5]), .QN());
   DFF_X1 \mem_reg[13][4]  (.D(n_0_612), .CK(n_0), .Q(\mem[13] [4]), .QN());
   DFF_X1 \mem_reg[13][3]  (.D(n_0_611), .CK(n_0), .Q(\mem[13] [3]), .QN());
   DFF_X1 \mem_reg[13][2]  (.D(n_0_610), .CK(n_0), .Q(\mem[13] [2]), .QN());
   DFF_X1 \mem_reg[13][1]  (.D(n_0_609), .CK(n_0), .Q(\mem[13] [1]), .QN());
   DFF_X1 \mem_reg[13][0]  (.D(n_0_608), .CK(n_0), .Q(\mem[13] [0]), .QN());
   DFF_X1 \mem_reg[14][15]  (.D(n_0_607), .CK(n_0), .Q(\mem[14] [15]), .QN());
   DFF_X1 \mem_reg[14][14]  (.D(n_0_606), .CK(n_0), .Q(\mem[14] [14]), .QN());
   DFF_X1 \mem_reg[14][13]  (.D(n_0_605), .CK(n_0), .Q(\mem[14] [13]), .QN());
   DFF_X1 \mem_reg[14][12]  (.D(n_0_604), .CK(n_0), .Q(\mem[14] [12]), .QN());
   DFF_X1 \mem_reg[14][11]  (.D(n_0_603), .CK(n_0), .Q(\mem[14] [11]), .QN());
   DFF_X1 \mem_reg[14][10]  (.D(n_0_602), .CK(n_0), .Q(\mem[14] [10]), .QN());
   DFF_X1 \mem_reg[14][9]  (.D(n_0_601), .CK(n_0), .Q(\mem[14] [9]), .QN());
   DFF_X1 \mem_reg[14][8]  (.D(n_0_600), .CK(n_0), .Q(\mem[14] [8]), .QN());
   DFF_X1 \mem_reg[14][7]  (.D(n_0_599), .CK(n_0), .Q(\mem[14] [7]), .QN());
   DFF_X1 \mem_reg[14][6]  (.D(n_0_598), .CK(n_0), .Q(\mem[14] [6]), .QN());
   DFF_X1 \mem_reg[14][5]  (.D(n_0_597), .CK(n_0), .Q(\mem[14] [5]), .QN());
   DFF_X1 \mem_reg[14][4]  (.D(n_0_596), .CK(n_0), .Q(\mem[14] [4]), .QN());
   DFF_X1 \mem_reg[14][3]  (.D(n_0_595), .CK(n_0), .Q(\mem[14] [3]), .QN());
   DFF_X1 \mem_reg[14][2]  (.D(n_0_594), .CK(n_0), .Q(\mem[14] [2]), .QN());
   DFF_X1 \mem_reg[14][1]  (.D(n_0_593), .CK(n_0), .Q(\mem[14] [1]), .QN());
   DFF_X1 \mem_reg[14][0]  (.D(n_0_592), .CK(n_0), .Q(\mem[14] [0]), .QN());
   DFF_X1 \mem_reg[15][15]  (.D(n_0_591), .CK(n_0), .Q(\mem[15] [15]), .QN());
   DFF_X1 \mem_reg[15][14]  (.D(n_0_590), .CK(n_0), .Q(\mem[15] [14]), .QN());
   DFF_X1 \mem_reg[15][13]  (.D(n_0_589), .CK(n_0), .Q(\mem[15] [13]), .QN());
   DFF_X1 \mem_reg[15][12]  (.D(n_0_588), .CK(n_0), .Q(\mem[15] [12]), .QN());
   DFF_X1 \mem_reg[15][11]  (.D(n_0_587), .CK(n_0), .Q(\mem[15] [11]), .QN());
   DFF_X1 \mem_reg[15][10]  (.D(n_0_586), .CK(n_0), .Q(\mem[15] [10]), .QN());
   DFF_X1 \mem_reg[15][9]  (.D(n_0_585), .CK(n_0), .Q(\mem[15] [9]), .QN());
   DFF_X1 \mem_reg[15][8]  (.D(n_0_584), .CK(n_0), .Q(\mem[15] [8]), .QN());
   DFF_X1 \mem_reg[15][7]  (.D(n_0_583), .CK(n_0), .Q(\mem[15] [7]), .QN());
   DFF_X1 \mem_reg[15][6]  (.D(n_0_582), .CK(n_0), .Q(\mem[15] [6]), .QN());
   DFF_X1 \mem_reg[15][5]  (.D(n_0_581), .CK(n_0), .Q(\mem[15] [5]), .QN());
   DFF_X1 \mem_reg[15][4]  (.D(n_0_580), .CK(n_0), .Q(\mem[15] [4]), .QN());
   DFF_X1 \mem_reg[15][3]  (.D(n_0_579), .CK(n_0), .Q(\mem[15] [3]), .QN());
   DFF_X1 \mem_reg[15][2]  (.D(n_0_578), .CK(n_0), .Q(\mem[15] [2]), .QN());
   DFF_X1 \mem_reg[15][1]  (.D(n_0_577), .CK(n_0), .Q(\mem[15] [1]), .QN());
   DFF_X1 \mem_reg[15][0]  (.D(n_0_576), .CK(n_0), .Q(\mem[15] [0]), .QN());
   DFF_X1 \mem_reg[16][15]  (.D(n_0_575), .CK(n_0), .Q(\mem[16] [15]), .QN());
   DFF_X1 \mem_reg[16][14]  (.D(n_0_574), .CK(n_0), .Q(\mem[16] [14]), .QN());
   DFF_X1 \mem_reg[16][13]  (.D(n_0_573), .CK(n_0), .Q(\mem[16] [13]), .QN());
   DFF_X1 \mem_reg[16][12]  (.D(n_0_572), .CK(n_0), .Q(\mem[16] [12]), .QN());
   DFF_X1 \mem_reg[16][11]  (.D(n_0_571), .CK(n_0), .Q(\mem[16] [11]), .QN());
   DFF_X1 \mem_reg[16][10]  (.D(n_0_570), .CK(n_0), .Q(\mem[16] [10]), .QN());
   DFF_X1 \mem_reg[16][9]  (.D(n_0_569), .CK(n_0), .Q(\mem[16] [9]), .QN());
   DFF_X1 \mem_reg[16][8]  (.D(n_0_568), .CK(n_0), .Q(\mem[16] [8]), .QN());
   DFF_X1 \mem_reg[16][7]  (.D(n_0_567), .CK(n_0), .Q(\mem[16] [7]), .QN());
   DFF_X1 \mem_reg[16][6]  (.D(n_0_566), .CK(n_0), .Q(\mem[16] [6]), .QN());
   DFF_X1 \mem_reg[16][5]  (.D(n_0_565), .CK(n_0), .Q(\mem[16] [5]), .QN());
   DFF_X1 \mem_reg[16][4]  (.D(n_0_564), .CK(n_0), .Q(\mem[16] [4]), .QN());
   DFF_X1 \mem_reg[16][3]  (.D(n_0_563), .CK(n_0), .Q(\mem[16] [3]), .QN());
   DFF_X1 \mem_reg[16][2]  (.D(n_0_562), .CK(n_0), .Q(\mem[16] [2]), .QN());
   DFF_X1 \mem_reg[16][1]  (.D(n_0_561), .CK(n_0), .Q(\mem[16] [1]), .QN());
   DFF_X1 \mem_reg[16][0]  (.D(n_0_560), .CK(n_0), .Q(\mem[16] [0]), .QN());
   DFF_X1 \mem_reg[17][15]  (.D(n_0_559), .CK(n_0), .Q(\mem[17] [15]), .QN());
   DFF_X1 \mem_reg[17][14]  (.D(n_0_558), .CK(n_0), .Q(\mem[17] [14]), .QN());
   DFF_X1 \mem_reg[17][13]  (.D(n_0_557), .CK(n_0), .Q(\mem[17] [13]), .QN());
   DFF_X1 \mem_reg[17][12]  (.D(n_0_556), .CK(n_0), .Q(\mem[17] [12]), .QN());
   DFF_X1 \mem_reg[17][11]  (.D(n_0_555), .CK(n_0), .Q(\mem[17] [11]), .QN());
   DFF_X1 \mem_reg[17][10]  (.D(n_0_554), .CK(n_0), .Q(\mem[17] [10]), .QN());
   DFF_X1 \mem_reg[17][9]  (.D(n_0_553), .CK(n_0), .Q(\mem[17] [9]), .QN());
   DFF_X1 \mem_reg[17][8]  (.D(n_0_552), .CK(n_0), .Q(\mem[17] [8]), .QN());
   DFF_X1 \mem_reg[17][7]  (.D(n_0_551), .CK(n_0), .Q(\mem[17] [7]), .QN());
   DFF_X1 \mem_reg[17][6]  (.D(n_0_550), .CK(n_0), .Q(\mem[17] [6]), .QN());
   DFF_X1 \mem_reg[17][5]  (.D(n_0_549), .CK(n_0), .Q(\mem[17] [5]), .QN());
   DFF_X1 \mem_reg[17][4]  (.D(n_0_548), .CK(n_0), .Q(\mem[17] [4]), .QN());
   DFF_X1 \mem_reg[17][3]  (.D(n_0_547), .CK(n_0), .Q(\mem[17] [3]), .QN());
   DFF_X1 \mem_reg[17][2]  (.D(n_0_546), .CK(n_0), .Q(\mem[17] [2]), .QN());
   DFF_X1 \mem_reg[17][1]  (.D(n_0_545), .CK(n_0), .Q(\mem[17] [1]), .QN());
   DFF_X1 \mem_reg[17][0]  (.D(n_0_544), .CK(n_0), .Q(\mem[17] [0]), .QN());
   DFF_X1 \mem_reg[18][15]  (.D(n_0_543), .CK(n_0), .Q(\mem[18] [15]), .QN());
   DFF_X1 \mem_reg[18][14]  (.D(n_0_542), .CK(n_0), .Q(\mem[18] [14]), .QN());
   DFF_X1 \mem_reg[18][13]  (.D(n_0_541), .CK(n_0), .Q(\mem[18] [13]), .QN());
   DFF_X1 \mem_reg[18][12]  (.D(n_0_540), .CK(n_0), .Q(\mem[18] [12]), .QN());
   DFF_X1 \mem_reg[18][11]  (.D(n_0_539), .CK(n_0), .Q(\mem[18] [11]), .QN());
   DFF_X1 \mem_reg[18][10]  (.D(n_0_538), .CK(n_0), .Q(\mem[18] [10]), .QN());
   DFF_X1 \mem_reg[18][9]  (.D(n_0_537), .CK(n_0), .Q(\mem[18] [9]), .QN());
   DFF_X1 \mem_reg[18][8]  (.D(n_0_536), .CK(n_0), .Q(\mem[18] [8]), .QN());
   DFF_X1 \mem_reg[18][7]  (.D(n_0_535), .CK(n_0), .Q(\mem[18] [7]), .QN());
   DFF_X1 \mem_reg[18][6]  (.D(n_0_534), .CK(n_0), .Q(\mem[18] [6]), .QN());
   DFF_X1 \mem_reg[18][5]  (.D(n_0_533), .CK(n_0), .Q(\mem[18] [5]), .QN());
   DFF_X1 \mem_reg[18][4]  (.D(n_0_532), .CK(n_0), .Q(\mem[18] [4]), .QN());
   DFF_X1 \mem_reg[18][3]  (.D(n_0_531), .CK(n_0), .Q(\mem[18] [3]), .QN());
   DFF_X1 \mem_reg[18][2]  (.D(n_0_530), .CK(n_0), .Q(\mem[18] [2]), .QN());
   DFF_X1 \mem_reg[18][1]  (.D(n_0_529), .CK(n_0), .Q(\mem[18] [1]), .QN());
   DFF_X1 \mem_reg[18][0]  (.D(n_0_528), .CK(n_0), .Q(\mem[18] [0]), .QN());
   DFF_X1 \mem_reg[19][15]  (.D(n_0_527), .CK(n_0), .Q(\mem[19] [15]), .QN());
   DFF_X1 \mem_reg[19][14]  (.D(n_0_526), .CK(n_0), .Q(\mem[19] [14]), .QN());
   DFF_X1 \mem_reg[19][13]  (.D(n_0_525), .CK(n_0), .Q(\mem[19] [13]), .QN());
   DFF_X1 \mem_reg[19][12]  (.D(n_0_524), .CK(n_0), .Q(\mem[19] [12]), .QN());
   DFF_X1 \mem_reg[19][11]  (.D(n_0_523), .CK(n_0), .Q(\mem[19] [11]), .QN());
   DFF_X1 \mem_reg[19][10]  (.D(n_0_522), .CK(n_0), .Q(\mem[19] [10]), .QN());
   DFF_X1 \mem_reg[19][9]  (.D(n_0_521), .CK(n_0), .Q(\mem[19] [9]), .QN());
   DFF_X1 \mem_reg[19][8]  (.D(n_0_520), .CK(n_0), .Q(\mem[19] [8]), .QN());
   DFF_X1 \mem_reg[19][7]  (.D(n_0_519), .CK(n_0), .Q(\mem[19] [7]), .QN());
   DFF_X1 \mem_reg[19][6]  (.D(n_0_518), .CK(n_0), .Q(\mem[19] [6]), .QN());
   DFF_X1 \mem_reg[19][5]  (.D(n_0_517), .CK(n_0), .Q(\mem[19] [5]), .QN());
   DFF_X1 \mem_reg[19][4]  (.D(n_0_516), .CK(n_0), .Q(\mem[19] [4]), .QN());
   DFF_X1 \mem_reg[19][3]  (.D(n_0_515), .CK(n_0), .Q(\mem[19] [3]), .QN());
   DFF_X1 \mem_reg[19][2]  (.D(n_0_514), .CK(n_0), .Q(\mem[19] [2]), .QN());
   DFF_X1 \mem_reg[19][1]  (.D(n_0_513), .CK(n_0), .Q(\mem[19] [1]), .QN());
   DFF_X1 \mem_reg[19][0]  (.D(n_0_512), .CK(n_0), .Q(\mem[19] [0]), .QN());
   DFF_X1 \mem_reg[20][15]  (.D(n_0_511), .CK(n_0), .Q(\mem[20] [15]), .QN());
   DFF_X1 \mem_reg[20][14]  (.D(n_0_510), .CK(n_0), .Q(\mem[20] [14]), .QN());
   DFF_X1 \mem_reg[20][13]  (.D(n_0_509), .CK(n_0), .Q(\mem[20] [13]), .QN());
   DFF_X1 \mem_reg[20][12]  (.D(n_0_508), .CK(n_0), .Q(\mem[20] [12]), .QN());
   DFF_X1 \mem_reg[20][11]  (.D(n_0_507), .CK(n_0), .Q(\mem[20] [11]), .QN());
   DFF_X1 \mem_reg[20][10]  (.D(n_0_506), .CK(n_0), .Q(\mem[20] [10]), .QN());
   DFF_X1 \mem_reg[20][9]  (.D(n_0_505), .CK(n_0), .Q(\mem[20] [9]), .QN());
   DFF_X1 \mem_reg[20][8]  (.D(n_0_504), .CK(n_0), .Q(\mem[20] [8]), .QN());
   DFF_X1 \mem_reg[20][7]  (.D(n_0_503), .CK(n_0), .Q(\mem[20] [7]), .QN());
   DFF_X1 \mem_reg[20][6]  (.D(n_0_502), .CK(n_0), .Q(\mem[20] [6]), .QN());
   DFF_X1 \mem_reg[20][5]  (.D(n_0_501), .CK(n_0), .Q(\mem[20] [5]), .QN());
   DFF_X1 \mem_reg[20][4]  (.D(n_0_500), .CK(n_0), .Q(\mem[20] [4]), .QN());
   DFF_X1 \mem_reg[20][3]  (.D(n_0_499), .CK(n_0), .Q(\mem[20] [3]), .QN());
   DFF_X1 \mem_reg[20][2]  (.D(n_0_498), .CK(n_0), .Q(\mem[20] [2]), .QN());
   DFF_X1 \mem_reg[20][1]  (.D(n_0_497), .CK(n_0), .Q(\mem[20] [1]), .QN());
   DFF_X1 \mem_reg[20][0]  (.D(n_0_496), .CK(n_0), .Q(\mem[20] [0]), .QN());
   DFF_X1 \mem_reg[21][15]  (.D(n_0_495), .CK(n_0), .Q(\mem[21] [15]), .QN());
   DFF_X1 \mem_reg[21][14]  (.D(n_0_494), .CK(n_0), .Q(\mem[21] [14]), .QN());
   DFF_X1 \mem_reg[21][13]  (.D(n_0_493), .CK(n_0), .Q(\mem[21] [13]), .QN());
   DFF_X1 \mem_reg[21][12]  (.D(n_0_492), .CK(n_0), .Q(\mem[21] [12]), .QN());
   DFF_X1 \mem_reg[21][11]  (.D(n_0_491), .CK(n_0), .Q(\mem[21] [11]), .QN());
   DFF_X1 \mem_reg[21][10]  (.D(n_0_490), .CK(n_0), .Q(\mem[21] [10]), .QN());
   DFF_X1 \mem_reg[21][9]  (.D(n_0_489), .CK(n_0), .Q(\mem[21] [9]), .QN());
   DFF_X1 \mem_reg[21][8]  (.D(n_0_488), .CK(n_0), .Q(\mem[21] [8]), .QN());
   DFF_X1 \mem_reg[21][7]  (.D(n_0_487), .CK(n_0), .Q(\mem[21] [7]), .QN());
   DFF_X1 \mem_reg[21][6]  (.D(n_0_486), .CK(n_0), .Q(\mem[21] [6]), .QN());
   DFF_X1 \mem_reg[21][5]  (.D(n_0_485), .CK(n_0), .Q(\mem[21] [5]), .QN());
   DFF_X1 \mem_reg[21][4]  (.D(n_0_484), .CK(n_0), .Q(\mem[21] [4]), .QN());
   DFF_X1 \mem_reg[21][3]  (.D(n_0_483), .CK(n_0), .Q(\mem[21] [3]), .QN());
   DFF_X1 \mem_reg[21][2]  (.D(n_0_482), .CK(n_0), .Q(\mem[21] [2]), .QN());
   DFF_X1 \mem_reg[21][1]  (.D(n_0_481), .CK(n_0), .Q(\mem[21] [1]), .QN());
   DFF_X1 \mem_reg[21][0]  (.D(n_0_480), .CK(n_0), .Q(\mem[21] [0]), .QN());
   DFF_X1 \mem_reg[22][15]  (.D(n_0_479), .CK(n_0), .Q(\mem[22] [15]), .QN());
   DFF_X1 \mem_reg[22][14]  (.D(n_0_478), .CK(n_0), .Q(\mem[22] [14]), .QN());
   DFF_X1 \mem_reg[22][13]  (.D(n_0_477), .CK(n_0), .Q(\mem[22] [13]), .QN());
   DFF_X1 \mem_reg[22][12]  (.D(n_0_476), .CK(n_0), .Q(\mem[22] [12]), .QN());
   DFF_X1 \mem_reg[22][11]  (.D(n_0_475), .CK(n_0), .Q(\mem[22] [11]), .QN());
   DFF_X1 \mem_reg[22][10]  (.D(n_0_474), .CK(n_0), .Q(\mem[22] [10]), .QN());
   DFF_X1 \mem_reg[22][9]  (.D(n_0_473), .CK(n_0), .Q(\mem[22] [9]), .QN());
   DFF_X1 \mem_reg[22][8]  (.D(n_0_472), .CK(n_0), .Q(\mem[22] [8]), .QN());
   DFF_X1 \mem_reg[22][7]  (.D(n_0_471), .CK(n_0), .Q(\mem[22] [7]), .QN());
   DFF_X1 \mem_reg[22][6]  (.D(n_0_470), .CK(n_0), .Q(\mem[22] [6]), .QN());
   DFF_X1 \mem_reg[22][5]  (.D(n_0_469), .CK(n_0), .Q(\mem[22] [5]), .QN());
   DFF_X1 \mem_reg[22][4]  (.D(n_0_468), .CK(n_0), .Q(\mem[22] [4]), .QN());
   DFF_X1 \mem_reg[22][3]  (.D(n_0_467), .CK(n_0), .Q(\mem[22] [3]), .QN());
   DFF_X1 \mem_reg[22][2]  (.D(n_0_466), .CK(n_0), .Q(\mem[22] [2]), .QN());
   DFF_X1 \mem_reg[22][1]  (.D(n_0_465), .CK(n_0), .Q(\mem[22] [1]), .QN());
   DFF_X1 \mem_reg[22][0]  (.D(n_0_464), .CK(n_0), .Q(\mem[22] [0]), .QN());
   DFF_X1 \mem_reg[23][15]  (.D(n_0_463), .CK(n_0), .Q(\mem[23] [15]), .QN());
   DFF_X1 \mem_reg[23][14]  (.D(n_0_462), .CK(n_0), .Q(\mem[23] [14]), .QN());
   DFF_X1 \mem_reg[23][13]  (.D(n_0_461), .CK(n_0), .Q(\mem[23] [13]), .QN());
   DFF_X1 \mem_reg[23][12]  (.D(n_0_460), .CK(n_0), .Q(\mem[23] [12]), .QN());
   DFF_X1 \mem_reg[23][11]  (.D(n_0_459), .CK(n_0), .Q(\mem[23] [11]), .QN());
   DFF_X1 \mem_reg[23][10]  (.D(n_0_458), .CK(n_0), .Q(\mem[23] [10]), .QN());
   DFF_X1 \mem_reg[23][9]  (.D(n_0_457), .CK(n_0), .Q(\mem[23] [9]), .QN());
   DFF_X1 \mem_reg[23][8]  (.D(n_0_456), .CK(n_0), .Q(\mem[23] [8]), .QN());
   DFF_X1 \mem_reg[23][7]  (.D(n_0_455), .CK(n_0), .Q(\mem[23] [7]), .QN());
   DFF_X1 \mem_reg[23][6]  (.D(n_0_454), .CK(n_0), .Q(\mem[23] [6]), .QN());
   DFF_X1 \mem_reg[23][5]  (.D(n_0_453), .CK(n_0), .Q(\mem[23] [5]), .QN());
   DFF_X1 \mem_reg[23][4]  (.D(n_0_452), .CK(n_0), .Q(\mem[23] [4]), .QN());
   DFF_X1 \mem_reg[23][3]  (.D(n_0_451), .CK(n_0), .Q(\mem[23] [3]), .QN());
   DFF_X1 \mem_reg[23][2]  (.D(n_0_450), .CK(n_0), .Q(\mem[23] [2]), .QN());
   DFF_X1 \mem_reg[23][1]  (.D(n_0_449), .CK(n_0), .Q(\mem[23] [1]), .QN());
   DFF_X1 \mem_reg[23][0]  (.D(n_0_448), .CK(n_0), .Q(\mem[23] [0]), .QN());
   DFF_X1 \mem_reg[24][15]  (.D(n_0_447), .CK(n_0), .Q(\mem[24] [15]), .QN());
   DFF_X1 \mem_reg[24][14]  (.D(n_0_446), .CK(n_0), .Q(\mem[24] [14]), .QN());
   DFF_X1 \mem_reg[24][13]  (.D(n_0_445), .CK(n_0), .Q(\mem[24] [13]), .QN());
   DFF_X1 \mem_reg[24][12]  (.D(n_0_444), .CK(n_0), .Q(\mem[24] [12]), .QN());
   DFF_X1 \mem_reg[24][11]  (.D(n_0_443), .CK(n_0), .Q(\mem[24] [11]), .QN());
   DFF_X1 \mem_reg[24][10]  (.D(n_0_442), .CK(n_0), .Q(\mem[24] [10]), .QN());
   DFF_X1 \mem_reg[24][9]  (.D(n_0_441), .CK(n_0), .Q(\mem[24] [9]), .QN());
   DFF_X1 \mem_reg[24][8]  (.D(n_0_440), .CK(n_0), .Q(\mem[24] [8]), .QN());
   DFF_X1 \mem_reg[24][7]  (.D(n_0_439), .CK(n_0), .Q(\mem[24] [7]), .QN());
   DFF_X1 \mem_reg[24][6]  (.D(n_0_438), .CK(n_0), .Q(\mem[24] [6]), .QN());
   DFF_X1 \mem_reg[24][5]  (.D(n_0_437), .CK(n_0), .Q(\mem[24] [5]), .QN());
   DFF_X1 \mem_reg[24][4]  (.D(n_0_436), .CK(n_0), .Q(\mem[24] [4]), .QN());
   DFF_X1 \mem_reg[24][3]  (.D(n_0_435), .CK(n_0), .Q(\mem[24] [3]), .QN());
   DFF_X1 \mem_reg[24][2]  (.D(n_0_434), .CK(n_0), .Q(\mem[24] [2]), .QN());
   DFF_X1 \mem_reg[24][1]  (.D(n_0_433), .CK(n_0), .Q(\mem[24] [1]), .QN());
   DFF_X1 \mem_reg[24][0]  (.D(n_0_432), .CK(n_0), .Q(\mem[24] [0]), .QN());
   DFF_X1 \mem_reg[25][15]  (.D(n_0_431), .CK(n_0), .Q(\mem[25] [15]), .QN());
   DFF_X1 \mem_reg[25][14]  (.D(n_0_430), .CK(n_0), .Q(\mem[25] [14]), .QN());
   DFF_X1 \mem_reg[25][13]  (.D(n_0_429), .CK(n_0), .Q(\mem[25] [13]), .QN());
   DFF_X1 \mem_reg[25][12]  (.D(n_0_428), .CK(n_0), .Q(\mem[25] [12]), .QN());
   DFF_X1 \mem_reg[25][11]  (.D(n_0_427), .CK(n_0), .Q(\mem[25] [11]), .QN());
   DFF_X1 \mem_reg[25][10]  (.D(n_0_426), .CK(n_0), .Q(\mem[25] [10]), .QN());
   DFF_X1 \mem_reg[25][9]  (.D(n_0_425), .CK(n_0), .Q(\mem[25] [9]), .QN());
   DFF_X1 \mem_reg[25][8]  (.D(n_0_424), .CK(n_0), .Q(\mem[25] [8]), .QN());
   DFF_X1 \mem_reg[25][7]  (.D(n_0_423), .CK(n_0), .Q(\mem[25] [7]), .QN());
   DFF_X1 \mem_reg[25][6]  (.D(n_0_422), .CK(n_0), .Q(\mem[25] [6]), .QN());
   DFF_X1 \mem_reg[25][5]  (.D(n_0_421), .CK(n_0), .Q(\mem[25] [5]), .QN());
   DFF_X1 \mem_reg[25][4]  (.D(n_0_420), .CK(n_0), .Q(\mem[25] [4]), .QN());
   DFF_X1 \mem_reg[25][3]  (.D(n_0_419), .CK(n_0), .Q(\mem[25] [3]), .QN());
   DFF_X1 \mem_reg[25][2]  (.D(n_0_418), .CK(n_0), .Q(\mem[25] [2]), .QN());
   DFF_X1 \mem_reg[25][1]  (.D(n_0_417), .CK(n_0), .Q(\mem[25] [1]), .QN());
   DFF_X1 \mem_reg[25][0]  (.D(n_0_416), .CK(n_0), .Q(\mem[25] [0]), .QN());
   DFF_X1 \mem_reg[26][15]  (.D(n_0_415), .CK(n_0), .Q(\mem[26] [15]), .QN());
   DFF_X1 \mem_reg[26][14]  (.D(n_0_414), .CK(n_0), .Q(\mem[26] [14]), .QN());
   DFF_X1 \mem_reg[26][13]  (.D(n_0_413), .CK(n_0), .Q(\mem[26] [13]), .QN());
   DFF_X1 \mem_reg[26][12]  (.D(n_0_412), .CK(n_0), .Q(\mem[26] [12]), .QN());
   DFF_X1 \mem_reg[26][11]  (.D(n_0_411), .CK(n_0), .Q(\mem[26] [11]), .QN());
   DFF_X1 \mem_reg[26][10]  (.D(n_0_410), .CK(n_0), .Q(\mem[26] [10]), .QN());
   DFF_X1 \mem_reg[26][9]  (.D(n_0_409), .CK(n_0), .Q(\mem[26] [9]), .QN());
   DFF_X1 \mem_reg[26][8]  (.D(n_0_408), .CK(n_0), .Q(\mem[26] [8]), .QN());
   DFF_X1 \mem_reg[26][7]  (.D(n_0_407), .CK(n_0), .Q(\mem[26] [7]), .QN());
   DFF_X1 \mem_reg[26][6]  (.D(n_0_406), .CK(n_0), .Q(\mem[26] [6]), .QN());
   DFF_X1 \mem_reg[26][5]  (.D(n_0_405), .CK(n_0), .Q(\mem[26] [5]), .QN());
   DFF_X1 \mem_reg[26][4]  (.D(n_0_404), .CK(n_0), .Q(\mem[26] [4]), .QN());
   DFF_X1 \mem_reg[26][3]  (.D(n_0_403), .CK(n_0), .Q(\mem[26] [3]), .QN());
   DFF_X1 \mem_reg[26][2]  (.D(n_0_402), .CK(n_0), .Q(\mem[26] [2]), .QN());
   DFF_X1 \mem_reg[26][1]  (.D(n_0_401), .CK(n_0), .Q(\mem[26] [1]), .QN());
   DFF_X1 \mem_reg[26][0]  (.D(n_0_400), .CK(n_0), .Q(\mem[26] [0]), .QN());
   DFF_X1 \mem_reg[27][15]  (.D(n_0_399), .CK(n_0), .Q(\mem[27] [15]), .QN());
   DFF_X1 \mem_reg[27][14]  (.D(n_0_398), .CK(n_0), .Q(\mem[27] [14]), .QN());
   DFF_X1 \mem_reg[27][13]  (.D(n_0_397), .CK(n_0), .Q(\mem[27] [13]), .QN());
   DFF_X1 \mem_reg[27][12]  (.D(n_0_396), .CK(n_0), .Q(\mem[27] [12]), .QN());
   DFF_X1 \mem_reg[27][11]  (.D(n_0_395), .CK(n_0), .Q(\mem[27] [11]), .QN());
   DFF_X1 \mem_reg[27][10]  (.D(n_0_394), .CK(n_0), .Q(\mem[27] [10]), .QN());
   DFF_X1 \mem_reg[27][9]  (.D(n_0_393), .CK(n_0), .Q(\mem[27] [9]), .QN());
   DFF_X1 \mem_reg[27][8]  (.D(n_0_392), .CK(n_0), .Q(\mem[27] [8]), .QN());
   DFF_X1 \mem_reg[27][7]  (.D(n_0_391), .CK(n_0), .Q(\mem[27] [7]), .QN());
   DFF_X1 \mem_reg[27][6]  (.D(n_0_390), .CK(n_0), .Q(\mem[27] [6]), .QN());
   DFF_X1 \mem_reg[27][5]  (.D(n_0_389), .CK(n_0), .Q(\mem[27] [5]), .QN());
   DFF_X1 \mem_reg[27][4]  (.D(n_0_388), .CK(n_0), .Q(\mem[27] [4]), .QN());
   DFF_X1 \mem_reg[27][3]  (.D(n_0_387), .CK(n_0), .Q(\mem[27] [3]), .QN());
   DFF_X1 \mem_reg[27][2]  (.D(n_0_386), .CK(n_0), .Q(\mem[27] [2]), .QN());
   DFF_X1 \mem_reg[27][1]  (.D(n_0_385), .CK(n_0), .Q(\mem[27] [1]), .QN());
   DFF_X1 \mem_reg[27][0]  (.D(n_0_384), .CK(n_0), .Q(\mem[27] [0]), .QN());
   DFF_X1 \mem_reg[28][15]  (.D(n_0_383), .CK(n_0), .Q(\mem[28] [15]), .QN());
   DFF_X1 \mem_reg[28][14]  (.D(n_0_382), .CK(n_0), .Q(\mem[28] [14]), .QN());
   DFF_X1 \mem_reg[28][13]  (.D(n_0_381), .CK(n_0), .Q(\mem[28] [13]), .QN());
   DFF_X1 \mem_reg[28][12]  (.D(n_0_380), .CK(n_0), .Q(\mem[28] [12]), .QN());
   DFF_X1 \mem_reg[28][11]  (.D(n_0_379), .CK(n_0), .Q(\mem[28] [11]), .QN());
   DFF_X1 \mem_reg[28][10]  (.D(n_0_378), .CK(n_0), .Q(\mem[28] [10]), .QN());
   DFF_X1 \mem_reg[28][9]  (.D(n_0_377), .CK(n_0), .Q(\mem[28] [9]), .QN());
   DFF_X1 \mem_reg[28][8]  (.D(n_0_376), .CK(n_0), .Q(\mem[28] [8]), .QN());
   DFF_X1 \mem_reg[28][7]  (.D(n_0_375), .CK(n_0), .Q(\mem[28] [7]), .QN());
   DFF_X1 \mem_reg[28][6]  (.D(n_0_374), .CK(n_0), .Q(\mem[28] [6]), .QN());
   DFF_X1 \mem_reg[28][5]  (.D(n_0_373), .CK(n_0), .Q(\mem[28] [5]), .QN());
   DFF_X1 \mem_reg[28][4]  (.D(n_0_372), .CK(n_0), .Q(\mem[28] [4]), .QN());
   DFF_X1 \mem_reg[28][3]  (.D(n_0_371), .CK(n_0), .Q(\mem[28] [3]), .QN());
   DFF_X1 \mem_reg[28][2]  (.D(n_0_370), .CK(n_0), .Q(\mem[28] [2]), .QN());
   DFF_X1 \mem_reg[28][1]  (.D(n_0_369), .CK(n_0), .Q(\mem[28] [1]), .QN());
   DFF_X1 \mem_reg[28][0]  (.D(n_0_368), .CK(n_0), .Q(\mem[28] [0]), .QN());
   DFF_X1 \mem_reg[29][15]  (.D(n_0_367), .CK(n_0), .Q(\mem[29] [15]), .QN());
   DFF_X1 \mem_reg[29][14]  (.D(n_0_366), .CK(n_0), .Q(\mem[29] [14]), .QN());
   DFF_X1 \mem_reg[29][13]  (.D(n_0_365), .CK(n_0), .Q(\mem[29] [13]), .QN());
   DFF_X1 \mem_reg[29][12]  (.D(n_0_364), .CK(n_0), .Q(\mem[29] [12]), .QN());
   DFF_X1 \mem_reg[29][11]  (.D(n_0_363), .CK(n_0), .Q(\mem[29] [11]), .QN());
   DFF_X1 \mem_reg[29][10]  (.D(n_0_362), .CK(n_0), .Q(\mem[29] [10]), .QN());
   DFF_X1 \mem_reg[29][9]  (.D(n_0_361), .CK(n_0), .Q(\mem[29] [9]), .QN());
   DFF_X1 \mem_reg[29][8]  (.D(n_0_360), .CK(n_0), .Q(\mem[29] [8]), .QN());
   DFF_X1 \mem_reg[29][7]  (.D(n_0_359), .CK(n_0), .Q(\mem[29] [7]), .QN());
   DFF_X1 \mem_reg[29][6]  (.D(n_0_358), .CK(n_0), .Q(\mem[29] [6]), .QN());
   DFF_X1 \mem_reg[29][5]  (.D(n_0_357), .CK(n_0), .Q(\mem[29] [5]), .QN());
   DFF_X1 \mem_reg[29][4]  (.D(n_0_356), .CK(n_0), .Q(\mem[29] [4]), .QN());
   DFF_X1 \mem_reg[29][3]  (.D(n_0_355), .CK(n_0), .Q(\mem[29] [3]), .QN());
   DFF_X1 \mem_reg[29][2]  (.D(n_0_354), .CK(n_0), .Q(\mem[29] [2]), .QN());
   DFF_X1 \mem_reg[29][1]  (.D(n_0_353), .CK(n_0), .Q(\mem[29] [1]), .QN());
   DFF_X1 \mem_reg[29][0]  (.D(n_0_352), .CK(n_0), .Q(\mem[29] [0]), .QN());
   DFF_X1 \mem_reg[30][15]  (.D(n_0_351), .CK(n_0), .Q(\mem[30] [15]), .QN());
   DFF_X1 \mem_reg[30][14]  (.D(n_0_350), .CK(n_0), .Q(\mem[30] [14]), .QN());
   DFF_X1 \mem_reg[30][13]  (.D(n_0_349), .CK(n_0), .Q(\mem[30] [13]), .QN());
   DFF_X1 \mem_reg[30][12]  (.D(n_0_348), .CK(n_0), .Q(\mem[30] [12]), .QN());
   DFF_X1 \mem_reg[30][11]  (.D(n_0_347), .CK(n_0), .Q(\mem[30] [11]), .QN());
   DFF_X1 \mem_reg[30][10]  (.D(n_0_346), .CK(n_0), .Q(\mem[30] [10]), .QN());
   DFF_X1 \mem_reg[30][9]  (.D(n_0_345), .CK(n_0), .Q(\mem[30] [9]), .QN());
   DFF_X1 \mem_reg[30][8]  (.D(n_0_344), .CK(n_0), .Q(\mem[30] [8]), .QN());
   DFF_X1 \mem_reg[30][7]  (.D(n_0_343), .CK(n_0), .Q(\mem[30] [7]), .QN());
   DFF_X1 \mem_reg[30][6]  (.D(n_0_342), .CK(n_0), .Q(\mem[30] [6]), .QN());
   DFF_X1 \mem_reg[30][5]  (.D(n_0_341), .CK(n_0), .Q(\mem[30] [5]), .QN());
   DFF_X1 \mem_reg[30][4]  (.D(n_0_340), .CK(n_0), .Q(\mem[30] [4]), .QN());
   DFF_X1 \mem_reg[30][3]  (.D(n_0_339), .CK(n_0), .Q(\mem[30] [3]), .QN());
   DFF_X1 \mem_reg[30][2]  (.D(n_0_338), .CK(n_0), .Q(\mem[30] [2]), .QN());
   DFF_X1 \mem_reg[30][1]  (.D(n_0_337), .CK(n_0), .Q(\mem[30] [1]), .QN());
   DFF_X1 \mem_reg[30][0]  (.D(n_0_336), .CK(n_0), .Q(\mem[30] [0]), .QN());
   DFF_X1 \mem_reg[31][15]  (.D(n_0_335), .CK(n_0), .Q(\mem[31] [15]), .QN());
   DFF_X1 \mem_reg[31][14]  (.D(n_0_334), .CK(n_0), .Q(\mem[31] [14]), .QN());
   DFF_X1 \mem_reg[31][13]  (.D(n_0_333), .CK(n_0), .Q(\mem[31] [13]), .QN());
   DFF_X1 \mem_reg[31][12]  (.D(n_0_332), .CK(n_0), .Q(\mem[31] [12]), .QN());
   DFF_X1 \mem_reg[31][11]  (.D(n_0_331), .CK(n_0), .Q(\mem[31] [11]), .QN());
   DFF_X1 \mem_reg[31][10]  (.D(n_0_330), .CK(n_0), .Q(\mem[31] [10]), .QN());
   DFF_X1 \mem_reg[31][9]  (.D(n_0_329), .CK(n_0), .Q(\mem[31] [9]), .QN());
   DFF_X1 \mem_reg[31][8]  (.D(n_0_328), .CK(n_0), .Q(\mem[31] [8]), .QN());
   DFF_X1 \mem_reg[31][7]  (.D(n_0_327), .CK(n_0), .Q(\mem[31] [7]), .QN());
   DFF_X1 \mem_reg[31][6]  (.D(n_0_326), .CK(n_0), .Q(\mem[31] [6]), .QN());
   DFF_X1 \mem_reg[31][5]  (.D(n_0_325), .CK(n_0), .Q(\mem[31] [5]), .QN());
   DFF_X1 \mem_reg[31][4]  (.D(n_0_324), .CK(n_0), .Q(\mem[31] [4]), .QN());
   DFF_X1 \mem_reg[31][3]  (.D(n_0_323), .CK(n_0), .Q(\mem[31] [3]), .QN());
   DFF_X1 \mem_reg[31][2]  (.D(n_0_322), .CK(n_0), .Q(\mem[31] [2]), .QN());
   DFF_X1 \mem_reg[31][1]  (.D(n_0_321), .CK(n_0), .Q(\mem[31] [1]), .QN());
   DFF_X1 \mem_reg[31][0]  (.D(n_0_320), .CK(n_0), .Q(\mem[31] [0]), .QN());
   DFF_X1 \mem_reg[32][15]  (.D(n_0_319), .CK(n_0), .Q(\mem[32] [15]), .QN());
   DFF_X1 \mem_reg[32][14]  (.D(n_0_318), .CK(n_0), .Q(\mem[32] [14]), .QN());
   DFF_X1 \mem_reg[32][13]  (.D(n_0_317), .CK(n_0), .Q(\mem[32] [13]), .QN());
   DFF_X1 \mem_reg[32][12]  (.D(n_0_316), .CK(n_0), .Q(\mem[32] [12]), .QN());
   DFF_X1 \mem_reg[32][11]  (.D(n_0_315), .CK(n_0), .Q(\mem[32] [11]), .QN());
   DFF_X1 \mem_reg[32][10]  (.D(n_0_314), .CK(n_0), .Q(\mem[32] [10]), .QN());
   DFF_X1 \mem_reg[32][9]  (.D(n_0_313), .CK(n_0), .Q(\mem[32] [9]), .QN());
   DFF_X1 \mem_reg[32][8]  (.D(n_0_312), .CK(n_0), .Q(\mem[32] [8]), .QN());
   DFF_X1 \mem_reg[32][7]  (.D(n_0_311), .CK(n_0), .Q(\mem[32] [7]), .QN());
   DFF_X1 \mem_reg[32][6]  (.D(n_0_310), .CK(n_0), .Q(\mem[32] [6]), .QN());
   DFF_X1 \mem_reg[32][5]  (.D(n_0_309), .CK(n_0), .Q(\mem[32] [5]), .QN());
   DFF_X1 \mem_reg[32][4]  (.D(n_0_308), .CK(n_0), .Q(\mem[32] [4]), .QN());
   DFF_X1 \mem_reg[32][3]  (.D(n_0_307), .CK(n_0), .Q(\mem[32] [3]), .QN());
   DFF_X1 \mem_reg[32][2]  (.D(n_0_306), .CK(n_0), .Q(\mem[32] [2]), .QN());
   DFF_X1 \mem_reg[32][1]  (.D(n_0_305), .CK(n_0), .Q(\mem[32] [1]), .QN());
   DFF_X1 \mem_reg[32][0]  (.D(n_0_304), .CK(n_0), .Q(\mem[32] [0]), .QN());
   DFF_X1 \mem_reg[33][15]  (.D(n_0_303), .CK(n_0), .Q(\mem[33] [15]), .QN());
   DFF_X1 \mem_reg[33][14]  (.D(n_0_302), .CK(n_0), .Q(\mem[33] [14]), .QN());
   DFF_X1 \mem_reg[33][13]  (.D(n_0_301), .CK(n_0), .Q(\mem[33] [13]), .QN());
   DFF_X1 \mem_reg[33][12]  (.D(n_0_300), .CK(n_0), .Q(\mem[33] [12]), .QN());
   DFF_X1 \mem_reg[33][11]  (.D(n_0_299), .CK(n_0), .Q(\mem[33] [11]), .QN());
   DFF_X1 \mem_reg[33][10]  (.D(n_0_298), .CK(n_0), .Q(\mem[33] [10]), .QN());
   DFF_X1 \mem_reg[33][9]  (.D(n_0_297), .CK(n_0), .Q(\mem[33] [9]), .QN());
   DFF_X1 \mem_reg[33][8]  (.D(n_0_296), .CK(n_0), .Q(\mem[33] [8]), .QN());
   DFF_X1 \mem_reg[33][7]  (.D(n_0_295), .CK(n_0), .Q(\mem[33] [7]), .QN());
   DFF_X1 \mem_reg[33][6]  (.D(n_0_294), .CK(n_0), .Q(\mem[33] [6]), .QN());
   DFF_X1 \mem_reg[33][5]  (.D(n_0_293), .CK(n_0), .Q(\mem[33] [5]), .QN());
   DFF_X1 \mem_reg[33][4]  (.D(n_0_292), .CK(n_0), .Q(\mem[33] [4]), .QN());
   DFF_X1 \mem_reg[33][3]  (.D(n_0_291), .CK(n_0), .Q(\mem[33] [3]), .QN());
   DFF_X1 \mem_reg[33][2]  (.D(n_0_290), .CK(n_0), .Q(\mem[33] [2]), .QN());
   DFF_X1 \mem_reg[33][1]  (.D(n_0_289), .CK(n_0), .Q(\mem[33] [1]), .QN());
   DFF_X1 \mem_reg[33][0]  (.D(n_0_288), .CK(n_0), .Q(\mem[33] [0]), .QN());
   DFF_X1 \mem_reg[34][15]  (.D(n_0_287), .CK(n_0), .Q(\mem[34] [15]), .QN());
   DFF_X1 \mem_reg[34][14]  (.D(n_0_286), .CK(n_0), .Q(\mem[34] [14]), .QN());
   DFF_X1 \mem_reg[34][13]  (.D(n_0_285), .CK(n_0), .Q(\mem[34] [13]), .QN());
   DFF_X1 \mem_reg[34][12]  (.D(n_0_284), .CK(n_0), .Q(\mem[34] [12]), .QN());
   DFF_X1 \mem_reg[34][11]  (.D(n_0_283), .CK(n_0), .Q(\mem[34] [11]), .QN());
   DFF_X1 \mem_reg[34][10]  (.D(n_0_282), .CK(n_0), .Q(\mem[34] [10]), .QN());
   DFF_X1 \mem_reg[34][9]  (.D(n_0_281), .CK(n_0), .Q(\mem[34] [9]), .QN());
   DFF_X1 \mem_reg[34][8]  (.D(n_0_280), .CK(n_0), .Q(\mem[34] [8]), .QN());
   DFF_X1 \mem_reg[34][7]  (.D(n_0_279), .CK(n_0), .Q(\mem[34] [7]), .QN());
   DFF_X1 \mem_reg[34][6]  (.D(n_0_278), .CK(n_0), .Q(\mem[34] [6]), .QN());
   DFF_X1 \mem_reg[34][5]  (.D(n_0_277), .CK(n_0), .Q(\mem[34] [5]), .QN());
   DFF_X1 \mem_reg[34][4]  (.D(n_0_276), .CK(n_0), .Q(\mem[34] [4]), .QN());
   DFF_X1 \mem_reg[34][3]  (.D(n_0_275), .CK(n_0), .Q(\mem[34] [3]), .QN());
   DFF_X1 \mem_reg[34][2]  (.D(n_0_274), .CK(n_0), .Q(\mem[34] [2]), .QN());
   DFF_X1 \mem_reg[34][1]  (.D(n_0_273), .CK(n_0), .Q(\mem[34] [1]), .QN());
   DFF_X1 \mem_reg[34][0]  (.D(n_0_272), .CK(n_0), .Q(\mem[34] [0]), .QN());
   DFF_X1 \mem_reg[35][15]  (.D(n_0_271), .CK(n_0), .Q(\mem[35] [15]), .QN());
   DFF_X1 \mem_reg[35][14]  (.D(n_0_270), .CK(n_0), .Q(\mem[35] [14]), .QN());
   DFF_X1 \mem_reg[35][13]  (.D(n_0_269), .CK(n_0), .Q(\mem[35] [13]), .QN());
   DFF_X1 \mem_reg[35][12]  (.D(n_0_268), .CK(n_0), .Q(\mem[35] [12]), .QN());
   DFF_X1 \mem_reg[35][11]  (.D(n_0_267), .CK(n_0), .Q(\mem[35] [11]), .QN());
   DFF_X1 \mem_reg[35][10]  (.D(n_0_266), .CK(n_0), .Q(\mem[35] [10]), .QN());
   DFF_X1 \mem_reg[35][9]  (.D(n_0_265), .CK(n_0), .Q(\mem[35] [9]), .QN());
   DFF_X1 \mem_reg[35][8]  (.D(n_0_264), .CK(n_0), .Q(\mem[35] [8]), .QN());
   DFF_X1 \mem_reg[35][7]  (.D(n_0_263), .CK(n_0), .Q(\mem[35] [7]), .QN());
   DFF_X1 \mem_reg[35][6]  (.D(n_0_262), .CK(n_0), .Q(\mem[35] [6]), .QN());
   DFF_X1 \mem_reg[35][5]  (.D(n_0_261), .CK(n_0), .Q(\mem[35] [5]), .QN());
   DFF_X1 \mem_reg[35][4]  (.D(n_0_260), .CK(n_0), .Q(\mem[35] [4]), .QN());
   DFF_X1 \mem_reg[35][3]  (.D(n_0_259), .CK(n_0), .Q(\mem[35] [3]), .QN());
   DFF_X1 \mem_reg[35][2]  (.D(n_0_258), .CK(n_0), .Q(\mem[35] [2]), .QN());
   DFF_X1 \mem_reg[35][1]  (.D(n_0_257), .CK(n_0), .Q(\mem[35] [1]), .QN());
   DFF_X1 \mem_reg[35][0]  (.D(n_0_256), .CK(n_0), .Q(\mem[35] [0]), .QN());
   DFF_X1 \mem_reg[36][15]  (.D(n_0_255), .CK(n_0), .Q(\mem[36] [15]), .QN());
   DFF_X1 \mem_reg[36][14]  (.D(n_0_254), .CK(n_0), .Q(\mem[36] [14]), .QN());
   DFF_X1 \mem_reg[36][13]  (.D(n_0_253), .CK(n_0), .Q(\mem[36] [13]), .QN());
   DFF_X1 \mem_reg[36][12]  (.D(n_0_252), .CK(n_0), .Q(\mem[36] [12]), .QN());
   DFF_X1 \mem_reg[36][11]  (.D(n_0_251), .CK(n_0), .Q(\mem[36] [11]), .QN());
   DFF_X1 \mem_reg[36][10]  (.D(n_0_250), .CK(n_0), .Q(\mem[36] [10]), .QN());
   DFF_X1 \mem_reg[36][9]  (.D(n_0_249), .CK(n_0), .Q(\mem[36] [9]), .QN());
   DFF_X1 \mem_reg[36][8]  (.D(n_0_248), .CK(n_0), .Q(\mem[36] [8]), .QN());
   DFF_X1 \mem_reg[36][7]  (.D(n_0_247), .CK(n_0), .Q(\mem[36] [7]), .QN());
   DFF_X1 \mem_reg[36][6]  (.D(n_0_246), .CK(n_0), .Q(\mem[36] [6]), .QN());
   DFF_X1 \mem_reg[36][5]  (.D(n_0_245), .CK(n_0), .Q(\mem[36] [5]), .QN());
   DFF_X1 \mem_reg[36][4]  (.D(n_0_244), .CK(n_0), .Q(\mem[36] [4]), .QN());
   DFF_X1 \mem_reg[36][3]  (.D(n_0_243), .CK(n_0), .Q(\mem[36] [3]), .QN());
   DFF_X1 \mem_reg[36][2]  (.D(n_0_242), .CK(n_0), .Q(\mem[36] [2]), .QN());
   DFF_X1 \mem_reg[36][1]  (.D(n_0_241), .CK(n_0), .Q(\mem[36] [1]), .QN());
   DFF_X1 \mem_reg[36][0]  (.D(n_0_240), .CK(n_0), .Q(\mem[36] [0]), .QN());
   DFF_X1 \mem_reg[37][15]  (.D(n_0_239), .CK(n_0), .Q(\mem[37] [15]), .QN());
   DFF_X1 \mem_reg[37][14]  (.D(n_0_238), .CK(n_0), .Q(\mem[37] [14]), .QN());
   DFF_X1 \mem_reg[37][13]  (.D(n_0_237), .CK(n_0), .Q(\mem[37] [13]), .QN());
   DFF_X1 \mem_reg[37][12]  (.D(n_0_236), .CK(n_0), .Q(\mem[37] [12]), .QN());
   DFF_X1 \mem_reg[37][11]  (.D(n_0_235), .CK(n_0), .Q(\mem[37] [11]), .QN());
   DFF_X1 \mem_reg[37][10]  (.D(n_0_234), .CK(n_0), .Q(\mem[37] [10]), .QN());
   DFF_X1 \mem_reg[37][9]  (.D(n_0_233), .CK(n_0), .Q(\mem[37] [9]), .QN());
   DFF_X1 \mem_reg[37][8]  (.D(n_0_232), .CK(n_0), .Q(\mem[37] [8]), .QN());
   DFF_X1 \mem_reg[37][7]  (.D(n_0_231), .CK(n_0), .Q(\mem[37] [7]), .QN());
   DFF_X1 \mem_reg[37][6]  (.D(n_0_230), .CK(n_0), .Q(\mem[37] [6]), .QN());
   DFF_X1 \mem_reg[37][5]  (.D(n_0_229), .CK(n_0), .Q(\mem[37] [5]), .QN());
   DFF_X1 \mem_reg[37][4]  (.D(n_0_228), .CK(n_0), .Q(\mem[37] [4]), .QN());
   DFF_X1 \mem_reg[37][3]  (.D(n_0_227), .CK(n_0), .Q(\mem[37] [3]), .QN());
   DFF_X1 \mem_reg[37][2]  (.D(n_0_226), .CK(n_0), .Q(\mem[37] [2]), .QN());
   DFF_X1 \mem_reg[37][1]  (.D(n_0_225), .CK(n_0), .Q(\mem[37] [1]), .QN());
   DFF_X1 \mem_reg[37][0]  (.D(n_0_224), .CK(n_0), .Q(\mem[37] [0]), .QN());
   DFF_X1 \mem_reg[38][15]  (.D(n_0_223), .CK(n_0), .Q(\mem[38] [15]), .QN());
   DFF_X1 \mem_reg[38][14]  (.D(n_0_222), .CK(n_0), .Q(\mem[38] [14]), .QN());
   DFF_X1 \mem_reg[38][13]  (.D(n_0_221), .CK(n_0), .Q(\mem[38] [13]), .QN());
   DFF_X1 \mem_reg[38][12]  (.D(n_0_220), .CK(n_0), .Q(\mem[38] [12]), .QN());
   DFF_X1 \mem_reg[38][11]  (.D(n_0_219), .CK(n_0), .Q(\mem[38] [11]), .QN());
   DFF_X1 \mem_reg[38][10]  (.D(n_0_218), .CK(n_0), .Q(\mem[38] [10]), .QN());
   DFF_X1 \mem_reg[38][9]  (.D(n_0_217), .CK(n_0), .Q(\mem[38] [9]), .QN());
   DFF_X1 \mem_reg[38][8]  (.D(n_0_216), .CK(n_0), .Q(\mem[38] [8]), .QN());
   DFF_X1 \mem_reg[38][7]  (.D(n_0_215), .CK(n_0), .Q(\mem[38] [7]), .QN());
   DFF_X1 \mem_reg[38][6]  (.D(n_0_214), .CK(n_0), .Q(\mem[38] [6]), .QN());
   DFF_X1 \mem_reg[38][5]  (.D(n_0_213), .CK(n_0), .Q(\mem[38] [5]), .QN());
   DFF_X1 \mem_reg[38][4]  (.D(n_0_212), .CK(n_0), .Q(\mem[38] [4]), .QN());
   DFF_X1 \mem_reg[38][3]  (.D(n_0_211), .CK(n_0), .Q(\mem[38] [3]), .QN());
   DFF_X1 \mem_reg[38][2]  (.D(n_0_210), .CK(n_0), .Q(\mem[38] [2]), .QN());
   DFF_X1 \mem_reg[38][1]  (.D(n_0_209), .CK(n_0), .Q(\mem[38] [1]), .QN());
   DFF_X1 \mem_reg[38][0]  (.D(n_0_208), .CK(n_0), .Q(\mem[38] [0]), .QN());
   DFF_X1 \mem_reg[39][15]  (.D(n_0_207), .CK(n_0), .Q(\mem[39] [15]), .QN());
   DFF_X1 \mem_reg[39][14]  (.D(n_0_206), .CK(n_0), .Q(\mem[39] [14]), .QN());
   DFF_X1 \mem_reg[39][13]  (.D(n_0_205), .CK(n_0), .Q(\mem[39] [13]), .QN());
   DFF_X1 \mem_reg[39][12]  (.D(n_0_204), .CK(n_0), .Q(\mem[39] [12]), .QN());
   DFF_X1 \mem_reg[39][11]  (.D(n_0_203), .CK(n_0), .Q(\mem[39] [11]), .QN());
   DFF_X1 \mem_reg[39][10]  (.D(n_0_202), .CK(n_0), .Q(\mem[39] [10]), .QN());
   DFF_X1 \mem_reg[39][9]  (.D(n_0_201), .CK(n_0), .Q(\mem[39] [9]), .QN());
   DFF_X1 \mem_reg[39][8]  (.D(n_0_200), .CK(n_0), .Q(\mem[39] [8]), .QN());
   DFF_X1 \mem_reg[39][7]  (.D(n_0_199), .CK(n_0), .Q(\mem[39] [7]), .QN());
   DFF_X1 \mem_reg[39][6]  (.D(n_0_198), .CK(n_0), .Q(\mem[39] [6]), .QN());
   DFF_X1 \mem_reg[39][5]  (.D(n_0_197), .CK(n_0), .Q(\mem[39] [5]), .QN());
   DFF_X1 \mem_reg[39][4]  (.D(n_0_196), .CK(n_0), .Q(\mem[39] [4]), .QN());
   DFF_X1 \mem_reg[39][3]  (.D(n_0_195), .CK(n_0), .Q(\mem[39] [3]), .QN());
   DFF_X1 \mem_reg[39][2]  (.D(n_0_194), .CK(n_0), .Q(\mem[39] [2]), .QN());
   DFF_X1 \mem_reg[39][1]  (.D(n_0_193), .CK(n_0), .Q(\mem[39] [1]), .QN());
   DFF_X1 \mem_reg[39][0]  (.D(n_0_192), .CK(n_0), .Q(\mem[39] [0]), .QN());
   DFF_X1 \mem_reg[40][15]  (.D(n_0_191), .CK(n_0), .Q(\mem[40] [15]), .QN());
   DFF_X1 \mem_reg[40][14]  (.D(n_0_190), .CK(n_0), .Q(\mem[40] [14]), .QN());
   DFF_X1 \mem_reg[40][13]  (.D(n_0_189), .CK(n_0), .Q(\mem[40] [13]), .QN());
   DFF_X1 \mem_reg[40][12]  (.D(n_0_188), .CK(n_0), .Q(\mem[40] [12]), .QN());
   DFF_X1 \mem_reg[40][11]  (.D(n_0_187), .CK(n_0), .Q(\mem[40] [11]), .QN());
   DFF_X1 \mem_reg[40][10]  (.D(n_0_186), .CK(n_0), .Q(\mem[40] [10]), .QN());
   DFF_X1 \mem_reg[40][9]  (.D(n_0_185), .CK(n_0), .Q(\mem[40] [9]), .QN());
   DFF_X1 \mem_reg[40][8]  (.D(n_0_184), .CK(n_0), .Q(\mem[40] [8]), .QN());
   DFF_X1 \mem_reg[40][7]  (.D(n_0_183), .CK(n_0), .Q(\mem[40] [7]), .QN());
   DFF_X1 \mem_reg[40][6]  (.D(n_0_182), .CK(n_0), .Q(\mem[40] [6]), .QN());
   DFF_X1 \mem_reg[40][5]  (.D(n_0_181), .CK(n_0), .Q(\mem[40] [5]), .QN());
   DFF_X1 \mem_reg[40][4]  (.D(n_0_180), .CK(n_0), .Q(\mem[40] [4]), .QN());
   DFF_X1 \mem_reg[40][3]  (.D(n_0_179), .CK(n_0), .Q(\mem[40] [3]), .QN());
   DFF_X1 \mem_reg[40][2]  (.D(n_0_178), .CK(n_0), .Q(\mem[40] [2]), .QN());
   DFF_X1 \mem_reg[40][1]  (.D(n_0_177), .CK(n_0), .Q(\mem[40] [1]), .QN());
   DFF_X1 \mem_reg[40][0]  (.D(n_0_176), .CK(n_0), .Q(\mem[40] [0]), .QN());
   DFF_X1 \mem_reg[41][15]  (.D(n_0_175), .CK(n_0), .Q(\mem[41] [15]), .QN());
   DFF_X1 \mem_reg[41][14]  (.D(n_0_174), .CK(n_0), .Q(\mem[41] [14]), .QN());
   DFF_X1 \mem_reg[41][13]  (.D(n_0_173), .CK(n_0), .Q(\mem[41] [13]), .QN());
   DFF_X1 \mem_reg[41][12]  (.D(n_0_172), .CK(n_0), .Q(\mem[41] [12]), .QN());
   DFF_X1 \mem_reg[41][11]  (.D(n_0_171), .CK(n_0), .Q(\mem[41] [11]), .QN());
   DFF_X1 \mem_reg[41][10]  (.D(n_0_170), .CK(n_0), .Q(\mem[41] [10]), .QN());
   DFF_X1 \mem_reg[41][9]  (.D(n_0_169), .CK(n_0), .Q(\mem[41] [9]), .QN());
   DFF_X1 \mem_reg[41][8]  (.D(n_0_168), .CK(n_0), .Q(\mem[41] [8]), .QN());
   DFF_X1 \mem_reg[41][7]  (.D(n_0_167), .CK(n_0), .Q(\mem[41] [7]), .QN());
   DFF_X1 \mem_reg[41][6]  (.D(n_0_166), .CK(n_0), .Q(\mem[41] [6]), .QN());
   DFF_X1 \mem_reg[41][5]  (.D(n_0_165), .CK(n_0), .Q(\mem[41] [5]), .QN());
   DFF_X1 \mem_reg[41][4]  (.D(n_0_164), .CK(n_0), .Q(\mem[41] [4]), .QN());
   DFF_X1 \mem_reg[41][3]  (.D(n_0_163), .CK(n_0), .Q(\mem[41] [3]), .QN());
   DFF_X1 \mem_reg[41][2]  (.D(n_0_162), .CK(n_0), .Q(\mem[41] [2]), .QN());
   DFF_X1 \mem_reg[41][1]  (.D(n_0_161), .CK(n_0), .Q(\mem[41] [1]), .QN());
   DFF_X1 \mem_reg[41][0]  (.D(n_0_160), .CK(n_0), .Q(\mem[41] [0]), .QN());
   DFF_X1 \mem_reg[42][15]  (.D(n_0_159), .CK(n_0), .Q(\mem[42] [15]), .QN());
   DFF_X1 \mem_reg[42][14]  (.D(n_0_158), .CK(n_0), .Q(\mem[42] [14]), .QN());
   DFF_X1 \mem_reg[42][13]  (.D(n_0_157), .CK(n_0), .Q(\mem[42] [13]), .QN());
   DFF_X1 \mem_reg[42][12]  (.D(n_0_156), .CK(n_0), .Q(\mem[42] [12]), .QN());
   DFF_X1 \mem_reg[42][11]  (.D(n_0_155), .CK(n_0), .Q(\mem[42] [11]), .QN());
   DFF_X1 \mem_reg[42][10]  (.D(n_0_154), .CK(n_0), .Q(\mem[42] [10]), .QN());
   DFF_X1 \mem_reg[42][9]  (.D(n_0_153), .CK(n_0), .Q(\mem[42] [9]), .QN());
   DFF_X1 \mem_reg[42][8]  (.D(n_0_152), .CK(n_0), .Q(\mem[42] [8]), .QN());
   DFF_X1 \mem_reg[42][7]  (.D(n_0_151), .CK(n_0), .Q(\mem[42] [7]), .QN());
   DFF_X1 \mem_reg[42][6]  (.D(n_0_150), .CK(n_0), .Q(\mem[42] [6]), .QN());
   DFF_X1 \mem_reg[42][5]  (.D(n_0_149), .CK(n_0), .Q(\mem[42] [5]), .QN());
   DFF_X1 \mem_reg[42][4]  (.D(n_0_148), .CK(n_0), .Q(\mem[42] [4]), .QN());
   DFF_X1 \mem_reg[42][3]  (.D(n_0_147), .CK(n_0), .Q(\mem[42] [3]), .QN());
   DFF_X1 \mem_reg[42][2]  (.D(n_0_146), .CK(n_0), .Q(\mem[42] [2]), .QN());
   DFF_X1 \mem_reg[42][1]  (.D(n_0_145), .CK(n_0), .Q(\mem[42] [1]), .QN());
   DFF_X1 \mem_reg[42][0]  (.D(n_0_144), .CK(n_0), .Q(\mem[42] [0]), .QN());
   DFF_X1 \mem_reg[43][15]  (.D(n_0_143), .CK(n_0), .Q(\mem[43] [15]), .QN());
   DFF_X1 \mem_reg[43][14]  (.D(n_0_142), .CK(n_0), .Q(\mem[43] [14]), .QN());
   DFF_X1 \mem_reg[43][13]  (.D(n_0_141), .CK(n_0), .Q(\mem[43] [13]), .QN());
   DFF_X1 \mem_reg[43][12]  (.D(n_0_140), .CK(n_0), .Q(\mem[43] [12]), .QN());
   DFF_X1 \mem_reg[43][11]  (.D(n_0_139), .CK(n_0), .Q(\mem[43] [11]), .QN());
   DFF_X1 \mem_reg[43][10]  (.D(n_0_138), .CK(n_0), .Q(\mem[43] [10]), .QN());
   DFF_X1 \mem_reg[43][9]  (.D(n_0_137), .CK(n_0), .Q(\mem[43] [9]), .QN());
   DFF_X1 \mem_reg[43][8]  (.D(n_0_136), .CK(n_0), .Q(\mem[43] [8]), .QN());
   DFF_X1 \mem_reg[43][7]  (.D(n_0_135), .CK(n_0), .Q(\mem[43] [7]), .QN());
   DFF_X1 \mem_reg[43][6]  (.D(n_0_134), .CK(n_0), .Q(\mem[43] [6]), .QN());
   DFF_X1 \mem_reg[43][5]  (.D(n_0_133), .CK(n_0), .Q(\mem[43] [5]), .QN());
   DFF_X1 \mem_reg[43][4]  (.D(n_0_132), .CK(n_0), .Q(\mem[43] [4]), .QN());
   DFF_X1 \mem_reg[43][3]  (.D(n_0_131), .CK(n_0), .Q(\mem[43] [3]), .QN());
   DFF_X1 \mem_reg[43][2]  (.D(n_0_130), .CK(n_0), .Q(\mem[43] [2]), .QN());
   DFF_X1 \mem_reg[43][1]  (.D(n_0_129), .CK(n_0), .Q(\mem[43] [1]), .QN());
   DFF_X1 \mem_reg[43][0]  (.D(n_0_128), .CK(n_0), .Q(\mem[43] [0]), .QN());
   DFF_X1 \mem_reg[44][15]  (.D(n_0_127), .CK(n_0), .Q(\mem[44] [15]), .QN());
   DFF_X1 \mem_reg[44][14]  (.D(n_0_126), .CK(n_0), .Q(\mem[44] [14]), .QN());
   DFF_X1 \mem_reg[44][13]  (.D(n_0_125), .CK(n_0), .Q(\mem[44] [13]), .QN());
   DFF_X1 \mem_reg[44][12]  (.D(n_0_124), .CK(n_0), .Q(\mem[44] [12]), .QN());
   DFF_X1 \mem_reg[44][11]  (.D(n_0_123), .CK(n_0), .Q(\mem[44] [11]), .QN());
   DFF_X1 \mem_reg[44][10]  (.D(n_0_122), .CK(n_0), .Q(\mem[44] [10]), .QN());
   DFF_X1 \mem_reg[44][9]  (.D(n_0_121), .CK(n_0), .Q(\mem[44] [9]), .QN());
   DFF_X1 \mem_reg[44][8]  (.D(n_0_120), .CK(n_0), .Q(\mem[44] [8]), .QN());
   DFF_X1 \mem_reg[44][7]  (.D(n_0_119), .CK(n_0), .Q(\mem[44] [7]), .QN());
   DFF_X1 \mem_reg[44][6]  (.D(n_0_118), .CK(n_0), .Q(\mem[44] [6]), .QN());
   DFF_X1 \mem_reg[44][5]  (.D(n_0_117), .CK(n_0), .Q(\mem[44] [5]), .QN());
   DFF_X1 \mem_reg[44][4]  (.D(n_0_116), .CK(n_0), .Q(\mem[44] [4]), .QN());
   DFF_X1 \mem_reg[44][3]  (.D(n_0_115), .CK(n_0), .Q(\mem[44] [3]), .QN());
   DFF_X1 \mem_reg[44][2]  (.D(n_0_114), .CK(n_0), .Q(\mem[44] [2]), .QN());
   DFF_X1 \mem_reg[44][1]  (.D(n_0_113), .CK(n_0), .Q(\mem[44] [1]), .QN());
   DFF_X1 \mem_reg[44][0]  (.D(n_0_112), .CK(n_0), .Q(\mem[44] [0]), .QN());
   DFF_X1 \mem_reg[45][15]  (.D(n_0_111), .CK(n_0), .Q(\mem[45] [15]), .QN());
   DFF_X1 \mem_reg[45][14]  (.D(n_0_110), .CK(n_0), .Q(\mem[45] [14]), .QN());
   DFF_X1 \mem_reg[45][13]  (.D(n_0_109), .CK(n_0), .Q(\mem[45] [13]), .QN());
   DFF_X1 \mem_reg[45][12]  (.D(n_0_108), .CK(n_0), .Q(\mem[45] [12]), .QN());
   DFF_X1 \mem_reg[45][11]  (.D(n_0_107), .CK(n_0), .Q(\mem[45] [11]), .QN());
   DFF_X1 \mem_reg[45][10]  (.D(n_0_106), .CK(n_0), .Q(\mem[45] [10]), .QN());
   DFF_X1 \mem_reg[45][9]  (.D(n_0_105), .CK(n_0), .Q(\mem[45] [9]), .QN());
   DFF_X1 \mem_reg[45][8]  (.D(n_0_104), .CK(n_0), .Q(\mem[45] [8]), .QN());
   DFF_X1 \mem_reg[45][7]  (.D(n_0_103), .CK(n_0), .Q(\mem[45] [7]), .QN());
   DFF_X1 \mem_reg[45][6]  (.D(n_0_102), .CK(n_0), .Q(\mem[45] [6]), .QN());
   DFF_X1 \mem_reg[45][5]  (.D(n_0_101), .CK(n_0), .Q(\mem[45] [5]), .QN());
   DFF_X1 \mem_reg[45][4]  (.D(n_0_100), .CK(n_0), .Q(\mem[45] [4]), .QN());
   DFF_X1 \mem_reg[45][3]  (.D(n_0_99), .CK(n_0), .Q(\mem[45] [3]), .QN());
   DFF_X1 \mem_reg[45][2]  (.D(n_0_98), .CK(n_0), .Q(\mem[45] [2]), .QN());
   DFF_X1 \mem_reg[45][1]  (.D(n_0_97), .CK(n_0), .Q(\mem[45] [1]), .QN());
   DFF_X1 \mem_reg[45][0]  (.D(n_0_96), .CK(n_0), .Q(\mem[45] [0]), .QN());
   DFF_X1 \mem_reg[46][15]  (.D(n_0_95), .CK(n_0), .Q(\mem[46] [15]), .QN());
   DFF_X1 \mem_reg[46][14]  (.D(n_0_94), .CK(n_0), .Q(\mem[46] [14]), .QN());
   DFF_X1 \mem_reg[46][13]  (.D(n_0_93), .CK(n_0), .Q(\mem[46] [13]), .QN());
   DFF_X1 \mem_reg[46][12]  (.D(n_0_92), .CK(n_0), .Q(\mem[46] [12]), .QN());
   DFF_X1 \mem_reg[46][11]  (.D(n_0_91), .CK(n_0), .Q(\mem[46] [11]), .QN());
   DFF_X1 \mem_reg[46][10]  (.D(n_0_90), .CK(n_0), .Q(\mem[46] [10]), .QN());
   DFF_X1 \mem_reg[46][9]  (.D(n_0_89), .CK(n_0), .Q(\mem[46] [9]), .QN());
   DFF_X1 \mem_reg[46][8]  (.D(n_0_88), .CK(n_0), .Q(\mem[46] [8]), .QN());
   DFF_X1 \mem_reg[46][7]  (.D(n_0_87), .CK(n_0), .Q(\mem[46] [7]), .QN());
   DFF_X1 \mem_reg[46][6]  (.D(n_0_86), .CK(n_0), .Q(\mem[46] [6]), .QN());
   DFF_X1 \mem_reg[46][5]  (.D(n_0_85), .CK(n_0), .Q(\mem[46] [5]), .QN());
   DFF_X1 \mem_reg[46][4]  (.D(n_0_84), .CK(n_0), .Q(\mem[46] [4]), .QN());
   DFF_X1 \mem_reg[46][3]  (.D(n_0_83), .CK(n_0), .Q(\mem[46] [3]), .QN());
   DFF_X1 \mem_reg[46][2]  (.D(n_0_82), .CK(n_0), .Q(\mem[46] [2]), .QN());
   DFF_X1 \mem_reg[46][1]  (.D(n_0_81), .CK(n_0), .Q(\mem[46] [1]), .QN());
   DFF_X1 \mem_reg[46][0]  (.D(n_0_80), .CK(n_0), .Q(\mem[46] [0]), .QN());
   DFF_X1 \mem_reg[47][15]  (.D(n_0_79), .CK(n_0), .Q(\mem[47] [15]), .QN());
   DFF_X1 \mem_reg[47][14]  (.D(n_0_78), .CK(n_0), .Q(\mem[47] [14]), .QN());
   DFF_X1 \mem_reg[47][13]  (.D(n_0_77), .CK(n_0), .Q(\mem[47] [13]), .QN());
   DFF_X1 \mem_reg[47][12]  (.D(n_0_76), .CK(n_0), .Q(\mem[47] [12]), .QN());
   DFF_X1 \mem_reg[47][11]  (.D(n_0_75), .CK(n_0), .Q(\mem[47] [11]), .QN());
   DFF_X1 \mem_reg[47][10]  (.D(n_0_74), .CK(n_0), .Q(\mem[47] [10]), .QN());
   DFF_X1 \mem_reg[47][9]  (.D(n_0_73), .CK(n_0), .Q(\mem[47] [9]), .QN());
   DFF_X1 \mem_reg[47][8]  (.D(n_0_72), .CK(n_0), .Q(\mem[47] [8]), .QN());
   DFF_X1 \mem_reg[47][7]  (.D(n_0_71), .CK(n_0), .Q(\mem[47] [7]), .QN());
   DFF_X1 \mem_reg[47][6]  (.D(n_0_70), .CK(n_0), .Q(\mem[47] [6]), .QN());
   DFF_X1 \mem_reg[47][5]  (.D(n_0_69), .CK(n_0), .Q(\mem[47] [5]), .QN());
   DFF_X1 \mem_reg[47][4]  (.D(n_0_68), .CK(n_0), .Q(\mem[47] [4]), .QN());
   DFF_X1 \mem_reg[47][3]  (.D(n_0_67), .CK(n_0), .Q(\mem[47] [3]), .QN());
   DFF_X1 \mem_reg[47][2]  (.D(n_0_66), .CK(n_0), .Q(\mem[47] [2]), .QN());
   DFF_X1 \mem_reg[47][1]  (.D(n_0_65), .CK(n_0), .Q(\mem[47] [1]), .QN());
   DFF_X1 \mem_reg[47][0]  (.D(n_0_64), .CK(n_0), .Q(\mem[47] [0]), .QN());
   DFF_X1 \mem_reg[48][15]  (.D(n_0_63), .CK(n_0), .Q(\mem[48] [15]), .QN());
   DFF_X1 \mem_reg[48][14]  (.D(n_0_62), .CK(n_0), .Q(\mem[48] [14]), .QN());
   DFF_X1 \mem_reg[48][13]  (.D(n_0_61), .CK(n_0), .Q(\mem[48] [13]), .QN());
   DFF_X1 \mem_reg[48][12]  (.D(n_0_60), .CK(n_0), .Q(\mem[48] [12]), .QN());
   DFF_X1 \mem_reg[48][11]  (.D(n_0_59), .CK(n_0), .Q(\mem[48] [11]), .QN());
   DFF_X1 \mem_reg[48][10]  (.D(n_0_58), .CK(n_0), .Q(\mem[48] [10]), .QN());
   DFF_X1 \mem_reg[48][9]  (.D(n_0_57), .CK(n_0), .Q(\mem[48] [9]), .QN());
   DFF_X1 \mem_reg[48][8]  (.D(n_0_56), .CK(n_0), .Q(\mem[48] [8]), .QN());
   DFF_X1 \mem_reg[48][7]  (.D(n_0_55), .CK(n_0), .Q(\mem[48] [7]), .QN());
   DFF_X1 \mem_reg[48][6]  (.D(n_0_54), .CK(n_0), .Q(\mem[48] [6]), .QN());
   DFF_X1 \mem_reg[48][5]  (.D(n_0_53), .CK(n_0), .Q(\mem[48] [5]), .QN());
   DFF_X1 \mem_reg[48][4]  (.D(n_0_52), .CK(n_0), .Q(\mem[48] [4]), .QN());
   DFF_X1 \mem_reg[48][3]  (.D(n_0_51), .CK(n_0), .Q(\mem[48] [3]), .QN());
   DFF_X1 \mem_reg[48][2]  (.D(n_0_50), .CK(n_0), .Q(\mem[48] [2]), .QN());
   DFF_X1 \mem_reg[48][1]  (.D(n_0_49), .CK(n_0), .Q(\mem[48] [1]), .QN());
   DFF_X1 \mem_reg[48][0]  (.D(n_0_48), .CK(n_0), .Q(\mem[48] [0]), .QN());
   DFF_X1 \mem_reg[49][15]  (.D(n_0_47), .CK(n_0), .Q(\mem[49] [15]), .QN());
   DFF_X1 \mem_reg[49][14]  (.D(n_0_46), .CK(n_0), .Q(\mem[49] [14]), .QN());
   DFF_X1 \mem_reg[49][13]  (.D(n_0_45), .CK(n_0), .Q(\mem[49] [13]), .QN());
   DFF_X1 \mem_reg[49][12]  (.D(n_0_44), .CK(n_0), .Q(\mem[49] [12]), .QN());
   DFF_X1 \mem_reg[49][11]  (.D(n_0_43), .CK(n_0), .Q(\mem[49] [11]), .QN());
   DFF_X1 \mem_reg[49][10]  (.D(n_0_42), .CK(n_0), .Q(\mem[49] [10]), .QN());
   DFF_X1 \mem_reg[49][9]  (.D(n_0_41), .CK(n_0), .Q(\mem[49] [9]), .QN());
   DFF_X1 \mem_reg[49][8]  (.D(n_0_40), .CK(n_0), .Q(\mem[49] [8]), .QN());
   DFF_X1 \mem_reg[49][7]  (.D(n_0_39), .CK(n_0), .Q(\mem[49] [7]), .QN());
   DFF_X1 \mem_reg[49][6]  (.D(n_0_38), .CK(n_0), .Q(\mem[49] [6]), .QN());
   DFF_X1 \mem_reg[49][5]  (.D(n_0_37), .CK(n_0), .Q(\mem[49] [5]), .QN());
   DFF_X1 \mem_reg[49][4]  (.D(n_0_36), .CK(n_0), .Q(\mem[49] [4]), .QN());
   DFF_X1 \mem_reg[49][3]  (.D(n_0_35), .CK(n_0), .Q(\mem[49] [3]), .QN());
   DFF_X1 \mem_reg[49][2]  (.D(n_0_34), .CK(n_0), .Q(\mem[49] [2]), .QN());
   DFF_X1 \mem_reg[49][1]  (.D(n_0_33), .CK(n_0), .Q(\mem[49] [1]), .QN());
   DFF_X1 \mem_reg[49][0]  (.D(n_0_32), .CK(n_0), .Q(\mem[49] [0]), .QN());
   DFF_X1 \mem_reg[51][15]  (.D(n_0_31), .CK(n_0), .Q(\mem[51] [15]), .QN());
   DFF_X1 \mem_reg[51][14]  (.D(n_0_30), .CK(n_0), .Q(\mem[51] [14]), .QN());
   DFF_X1 \mem_reg[51][13]  (.D(n_0_29), .CK(n_0), .Q(\mem[51] [13]), .QN());
   DFF_X1 \mem_reg[51][12]  (.D(n_0_28), .CK(n_0), .Q(\mem[51] [12]), .QN());
   DFF_X1 \mem_reg[51][11]  (.D(n_0_27), .CK(n_0), .Q(\mem[51] [11]), .QN());
   DFF_X1 \mem_reg[51][10]  (.D(n_0_26), .CK(n_0), .Q(\mem[51] [10]), .QN());
   DFF_X1 \mem_reg[51][9]  (.D(n_0_25), .CK(n_0), .Q(\mem[51] [9]), .QN());
   DFF_X1 \mem_reg[51][8]  (.D(n_0_24), .CK(n_0), .Q(\mem[51] [8]), .QN());
   DFF_X1 \mem_reg[51][7]  (.D(n_0_23), .CK(n_0), .Q(\mem[51] [7]), .QN());
   DFF_X1 \mem_reg[51][6]  (.D(n_0_22), .CK(n_0), .Q(\mem[51] [6]), .QN());
   DFF_X1 \mem_reg[51][5]  (.D(n_0_21), .CK(n_0), .Q(\mem[51] [5]), .QN());
   DFF_X1 \mem_reg[51][4]  (.D(n_0_20), .CK(n_0), .Q(\mem[51] [4]), .QN());
   DFF_X1 \mem_reg[51][3]  (.D(n_0_19), .CK(n_0), .Q(\mem[51] [3]), .QN());
   DFF_X1 \mem_reg[51][2]  (.D(n_0_18), .CK(n_0), .Q(\mem[51] [2]), .QN());
   DFF_X1 \mem_reg[51][1]  (.D(n_0_17), .CK(n_0), .Q(\mem[51] [1]), .QN());
   DFF_X1 \mem_reg[51][0]  (.D(n_0_16), .CK(n_0), .Q(\mem[51] [0]), .QN());
   DFF_X1 \mem_reg[50][15]  (.D(n_0_15), .CK(n_0), .Q(\mem[50] [15]), .QN());
   DFF_X1 \mem_reg[50][14]  (.D(n_0_14), .CK(n_0), .Q(\mem[50] [14]), .QN());
   DFF_X1 \mem_reg[50][13]  (.D(n_0_13), .CK(n_0), .Q(\mem[50] [13]), .QN());
   DFF_X1 \mem_reg[50][12]  (.D(n_0_12), .CK(n_0), .Q(\mem[50] [12]), .QN());
   DFF_X1 \mem_reg[50][11]  (.D(n_0_11), .CK(n_0), .Q(\mem[50] [11]), .QN());
   DFF_X1 \mem_reg[50][10]  (.D(n_0_10), .CK(n_0), .Q(\mem[50] [10]), .QN());
   DFF_X1 \mem_reg[50][9]  (.D(n_0_9), .CK(n_0), .Q(\mem[50] [9]), .QN());
   DFF_X1 \mem_reg[50][8]  (.D(n_0_8), .CK(n_0), .Q(\mem[50] [8]), .QN());
   DFF_X1 \mem_reg[50][7]  (.D(n_0_7), .CK(n_0), .Q(\mem[50] [7]), .QN());
   DFF_X1 \mem_reg[50][6]  (.D(n_0_6), .CK(n_0), .Q(\mem[50] [6]), .QN());
   DFF_X1 \mem_reg[50][5]  (.D(n_0_5), .CK(n_0), .Q(\mem[50] [5]), .QN());
   DFF_X1 \mem_reg[50][4]  (.D(n_0_4), .CK(n_0), .Q(\mem[50] [4]), .QN());
   DFF_X1 \mem_reg[50][3]  (.D(n_0_3), .CK(n_0), .Q(\mem[50] [3]), .QN());
   DFF_X1 \mem_reg[50][2]  (.D(n_0_2), .CK(n_0), .Q(\mem[50] [2]), .QN());
   DFF_X1 \mem_reg[50][1]  (.D(n_0_1), .CK(n_0), .Q(\mem[50] [1]), .QN());
   DFF_X1 \mem_reg[50][0]  (.D(n_0_0), .CK(n_0), .Q(\mem[50] [0]), .QN());
   MUX2_X1 i_0_0_0 (.A(\mem[1] [15]), .B(data[15]), .S(n_2), .Z(n_0_815));
   MUX2_X1 i_0_0_1 (.A(\mem[1] [14]), .B(data[14]), .S(n_2), .Z(n_0_814));
   MUX2_X1 i_0_0_2 (.A(\mem[1] [13]), .B(data[13]), .S(n_2), .Z(n_0_813));
   MUX2_X1 i_0_0_3 (.A(\mem[1] [12]), .B(data[12]), .S(n_2), .Z(n_0_812));
   MUX2_X1 i_0_0_4 (.A(\mem[1] [11]), .B(data[11]), .S(n_2), .Z(n_0_811));
   MUX2_X1 i_0_0_5 (.A(\mem[1] [10]), .B(data[10]), .S(n_2), .Z(n_0_810));
   MUX2_X1 i_0_0_6 (.A(\mem[1] [9]), .B(data[9]), .S(n_2), .Z(n_0_809));
   MUX2_X1 i_0_0_7 (.A(\mem[1] [8]), .B(data[8]), .S(n_2), .Z(n_0_808));
   MUX2_X1 i_0_0_8 (.A(\mem[1] [7]), .B(data[7]), .S(n_2), .Z(n_0_807));
   MUX2_X1 i_0_0_9 (.A(\mem[1] [6]), .B(data[6]), .S(n_2), .Z(n_0_806));
   MUX2_X1 i_0_0_10 (.A(\mem[1] [5]), .B(data[5]), .S(n_2), .Z(n_0_805));
   MUX2_X1 i_0_0_11 (.A(\mem[1] [4]), .B(data[4]), .S(n_2), .Z(n_0_804));
   MUX2_X1 i_0_0_12 (.A(\mem[1] [3]), .B(data[3]), .S(n_2), .Z(n_0_803));
   MUX2_X1 i_0_0_13 (.A(\mem[1] [2]), .B(data[2]), .S(n_2), .Z(n_0_802));
   MUX2_X1 i_0_0_14 (.A(\mem[1] [1]), .B(data[1]), .S(n_2), .Z(n_0_801));
   MUX2_X1 i_0_0_15 (.A(\mem[1] [0]), .B(data[0]), .S(n_2), .Z(n_0_800));
   MUX2_X1 i_0_0_16 (.A(\mem[2] [15]), .B(data[15]), .S(n_3), .Z(n_0_799));
   MUX2_X1 i_0_0_17 (.A(\mem[2] [14]), .B(data[14]), .S(n_3), .Z(n_0_798));
   MUX2_X1 i_0_0_18 (.A(\mem[2] [13]), .B(data[13]), .S(n_3), .Z(n_0_797));
   MUX2_X1 i_0_0_19 (.A(\mem[2] [12]), .B(data[12]), .S(n_3), .Z(n_0_796));
   MUX2_X1 i_0_0_20 (.A(\mem[2] [11]), .B(data[11]), .S(n_3), .Z(n_0_795));
   MUX2_X1 i_0_0_21 (.A(\mem[2] [10]), .B(data[10]), .S(n_3), .Z(n_0_794));
   MUX2_X1 i_0_0_22 (.A(\mem[2] [9]), .B(data[9]), .S(n_3), .Z(n_0_793));
   MUX2_X1 i_0_0_23 (.A(\mem[2] [8]), .B(data[8]), .S(n_3), .Z(n_0_792));
   MUX2_X1 i_0_0_24 (.A(\mem[2] [7]), .B(data[7]), .S(n_3), .Z(n_0_791));
   MUX2_X1 i_0_0_25 (.A(\mem[2] [6]), .B(data[6]), .S(n_3), .Z(n_0_790));
   MUX2_X1 i_0_0_26 (.A(\mem[2] [5]), .B(data[5]), .S(n_3), .Z(n_0_789));
   MUX2_X1 i_0_0_27 (.A(\mem[2] [4]), .B(data[4]), .S(n_3), .Z(n_0_788));
   MUX2_X1 i_0_0_28 (.A(\mem[2] [3]), .B(data[3]), .S(n_3), .Z(n_0_787));
   MUX2_X1 i_0_0_29 (.A(\mem[2] [2]), .B(data[2]), .S(n_3), .Z(n_0_786));
   MUX2_X1 i_0_0_30 (.A(\mem[2] [1]), .B(data[1]), .S(n_3), .Z(n_0_785));
   MUX2_X1 i_0_0_31 (.A(\mem[2] [0]), .B(data[0]), .S(n_3), .Z(n_0_784));
   MUX2_X1 i_0_0_32 (.A(\mem[3] [15]), .B(data[15]), .S(n_4), .Z(n_0_783));
   MUX2_X1 i_0_0_33 (.A(\mem[3] [14]), .B(data[14]), .S(n_4), .Z(n_0_782));
   MUX2_X1 i_0_0_34 (.A(\mem[3] [13]), .B(data[13]), .S(n_4), .Z(n_0_781));
   MUX2_X1 i_0_0_35 (.A(\mem[3] [12]), .B(data[12]), .S(n_4), .Z(n_0_780));
   MUX2_X1 i_0_0_36 (.A(\mem[3] [11]), .B(data[11]), .S(n_4), .Z(n_0_779));
   MUX2_X1 i_0_0_37 (.A(\mem[3] [10]), .B(data[10]), .S(n_4), .Z(n_0_778));
   MUX2_X1 i_0_0_38 (.A(\mem[3] [9]), .B(data[9]), .S(n_4), .Z(n_0_777));
   MUX2_X1 i_0_0_39 (.A(\mem[3] [8]), .B(data[8]), .S(n_4), .Z(n_0_776));
   MUX2_X1 i_0_0_40 (.A(\mem[3] [7]), .B(data[7]), .S(n_4), .Z(n_0_775));
   MUX2_X1 i_0_0_41 (.A(\mem[3] [6]), .B(data[6]), .S(n_4), .Z(n_0_774));
   MUX2_X1 i_0_0_42 (.A(\mem[3] [5]), .B(data[5]), .S(n_4), .Z(n_0_773));
   MUX2_X1 i_0_0_43 (.A(\mem[3] [4]), .B(data[4]), .S(n_4), .Z(n_0_772));
   MUX2_X1 i_0_0_44 (.A(\mem[3] [3]), .B(data[3]), .S(n_4), .Z(n_0_771));
   MUX2_X1 i_0_0_45 (.A(\mem[3] [2]), .B(data[2]), .S(n_4), .Z(n_0_770));
   MUX2_X1 i_0_0_46 (.A(\mem[3] [1]), .B(data[1]), .S(n_4), .Z(n_0_769));
   MUX2_X1 i_0_0_47 (.A(\mem[3] [0]), .B(data[0]), .S(n_4), .Z(n_0_768));
   MUX2_X1 i_0_0_48 (.A(\mem[4] [15]), .B(data[15]), .S(n_5), .Z(n_0_767));
   MUX2_X1 i_0_0_49 (.A(\mem[4] [14]), .B(data[14]), .S(n_5), .Z(n_0_766));
   MUX2_X1 i_0_0_50 (.A(\mem[4] [13]), .B(data[13]), .S(n_5), .Z(n_0_765));
   MUX2_X1 i_0_0_51 (.A(\mem[4] [12]), .B(data[12]), .S(n_5), .Z(n_0_764));
   MUX2_X1 i_0_0_52 (.A(\mem[4] [11]), .B(data[11]), .S(n_5), .Z(n_0_763));
   MUX2_X1 i_0_0_53 (.A(\mem[4] [10]), .B(data[10]), .S(n_5), .Z(n_0_762));
   MUX2_X1 i_0_0_54 (.A(\mem[4] [9]), .B(data[9]), .S(n_5), .Z(n_0_761));
   MUX2_X1 i_0_0_55 (.A(\mem[4] [8]), .B(data[8]), .S(n_5), .Z(n_0_760));
   MUX2_X1 i_0_0_56 (.A(\mem[4] [7]), .B(data[7]), .S(n_5), .Z(n_0_759));
   MUX2_X1 i_0_0_57 (.A(\mem[4] [6]), .B(data[6]), .S(n_5), .Z(n_0_758));
   MUX2_X1 i_0_0_58 (.A(\mem[4] [5]), .B(data[5]), .S(n_5), .Z(n_0_757));
   MUX2_X1 i_0_0_59 (.A(\mem[4] [4]), .B(data[4]), .S(n_5), .Z(n_0_756));
   MUX2_X1 i_0_0_60 (.A(\mem[4] [3]), .B(data[3]), .S(n_5), .Z(n_0_755));
   MUX2_X1 i_0_0_61 (.A(\mem[4] [2]), .B(data[2]), .S(n_5), .Z(n_0_754));
   MUX2_X1 i_0_0_62 (.A(\mem[4] [1]), .B(data[1]), .S(n_5), .Z(n_0_753));
   MUX2_X1 i_0_0_63 (.A(\mem[4] [0]), .B(data[0]), .S(n_5), .Z(n_0_752));
   MUX2_X1 i_0_0_64 (.A(\mem[5] [15]), .B(data[15]), .S(n_6), .Z(n_0_751));
   MUX2_X1 i_0_0_65 (.A(\mem[5] [14]), .B(data[14]), .S(n_6), .Z(n_0_750));
   MUX2_X1 i_0_0_66 (.A(\mem[5] [13]), .B(data[13]), .S(n_6), .Z(n_0_749));
   MUX2_X1 i_0_0_67 (.A(\mem[5] [12]), .B(data[12]), .S(n_6), .Z(n_0_748));
   MUX2_X1 i_0_0_68 (.A(\mem[5] [11]), .B(data[11]), .S(n_6), .Z(n_0_747));
   MUX2_X1 i_0_0_69 (.A(\mem[5] [10]), .B(data[10]), .S(n_6), .Z(n_0_746));
   MUX2_X1 i_0_0_70 (.A(\mem[5] [9]), .B(data[9]), .S(n_6), .Z(n_0_745));
   MUX2_X1 i_0_0_71 (.A(\mem[5] [8]), .B(data[8]), .S(n_6), .Z(n_0_744));
   MUX2_X1 i_0_0_72 (.A(\mem[5] [7]), .B(data[7]), .S(n_6), .Z(n_0_743));
   MUX2_X1 i_0_0_73 (.A(\mem[5] [6]), .B(data[6]), .S(n_6), .Z(n_0_742));
   MUX2_X1 i_0_0_74 (.A(\mem[5] [5]), .B(data[5]), .S(n_6), .Z(n_0_741));
   MUX2_X1 i_0_0_75 (.A(\mem[5] [4]), .B(data[4]), .S(n_6), .Z(n_0_740));
   MUX2_X1 i_0_0_76 (.A(\mem[5] [3]), .B(data[3]), .S(n_6), .Z(n_0_739));
   MUX2_X1 i_0_0_77 (.A(\mem[5] [2]), .B(data[2]), .S(n_6), .Z(n_0_738));
   MUX2_X1 i_0_0_78 (.A(\mem[5] [1]), .B(data[1]), .S(n_6), .Z(n_0_737));
   MUX2_X1 i_0_0_79 (.A(\mem[5] [0]), .B(data[0]), .S(n_6), .Z(n_0_736));
   MUX2_X1 i_0_0_80 (.A(\mem[6] [15]), .B(data[15]), .S(n_7), .Z(n_0_735));
   MUX2_X1 i_0_0_81 (.A(\mem[6] [14]), .B(data[14]), .S(n_7), .Z(n_0_734));
   MUX2_X1 i_0_0_82 (.A(\mem[6] [13]), .B(data[13]), .S(n_7), .Z(n_0_733));
   MUX2_X1 i_0_0_83 (.A(\mem[6] [12]), .B(data[12]), .S(n_7), .Z(n_0_732));
   MUX2_X1 i_0_0_84 (.A(\mem[6] [11]), .B(data[11]), .S(n_7), .Z(n_0_731));
   MUX2_X1 i_0_0_85 (.A(\mem[6] [10]), .B(data[10]), .S(n_7), .Z(n_0_730));
   MUX2_X1 i_0_0_86 (.A(\mem[6] [9]), .B(data[9]), .S(n_7), .Z(n_0_729));
   MUX2_X1 i_0_0_87 (.A(\mem[6] [8]), .B(data[8]), .S(n_7), .Z(n_0_728));
   MUX2_X1 i_0_0_88 (.A(\mem[6] [7]), .B(data[7]), .S(n_7), .Z(n_0_727));
   MUX2_X1 i_0_0_89 (.A(\mem[6] [6]), .B(data[6]), .S(n_7), .Z(n_0_726));
   MUX2_X1 i_0_0_90 (.A(\mem[6] [5]), .B(data[5]), .S(n_7), .Z(n_0_725));
   MUX2_X1 i_0_0_91 (.A(\mem[6] [4]), .B(data[4]), .S(n_7), .Z(n_0_724));
   MUX2_X1 i_0_0_92 (.A(\mem[6] [3]), .B(data[3]), .S(n_7), .Z(n_0_723));
   MUX2_X1 i_0_0_93 (.A(\mem[6] [2]), .B(data[2]), .S(n_7), .Z(n_0_722));
   MUX2_X1 i_0_0_94 (.A(\mem[6] [1]), .B(data[1]), .S(n_7), .Z(n_0_721));
   MUX2_X1 i_0_0_95 (.A(\mem[6] [0]), .B(data[0]), .S(n_7), .Z(n_0_720));
   MUX2_X1 i_0_0_96 (.A(\mem[7] [15]), .B(data[15]), .S(n_8), .Z(n_0_719));
   MUX2_X1 i_0_0_97 (.A(\mem[7] [14]), .B(data[14]), .S(n_8), .Z(n_0_718));
   MUX2_X1 i_0_0_98 (.A(\mem[7] [13]), .B(data[13]), .S(n_8), .Z(n_0_717));
   MUX2_X1 i_0_0_99 (.A(\mem[7] [12]), .B(data[12]), .S(n_8), .Z(n_0_716));
   MUX2_X1 i_0_0_100 (.A(\mem[7] [11]), .B(data[11]), .S(n_8), .Z(n_0_715));
   MUX2_X1 i_0_0_101 (.A(\mem[7] [10]), .B(data[10]), .S(n_8), .Z(n_0_714));
   MUX2_X1 i_0_0_102 (.A(\mem[7] [9]), .B(data[9]), .S(n_8), .Z(n_0_713));
   MUX2_X1 i_0_0_103 (.A(\mem[7] [8]), .B(data[8]), .S(n_8), .Z(n_0_712));
   MUX2_X1 i_0_0_104 (.A(\mem[7] [7]), .B(data[7]), .S(n_8), .Z(n_0_711));
   MUX2_X1 i_0_0_105 (.A(\mem[7] [6]), .B(data[6]), .S(n_8), .Z(n_0_710));
   MUX2_X1 i_0_0_106 (.A(\mem[7] [5]), .B(data[5]), .S(n_8), .Z(n_0_709));
   MUX2_X1 i_0_0_107 (.A(\mem[7] [4]), .B(data[4]), .S(n_8), .Z(n_0_708));
   MUX2_X1 i_0_0_108 (.A(\mem[7] [3]), .B(data[3]), .S(n_8), .Z(n_0_707));
   MUX2_X1 i_0_0_109 (.A(\mem[7] [2]), .B(data[2]), .S(n_8), .Z(n_0_706));
   MUX2_X1 i_0_0_110 (.A(\mem[7] [1]), .B(data[1]), .S(n_8), .Z(n_0_705));
   MUX2_X1 i_0_0_111 (.A(\mem[7] [0]), .B(data[0]), .S(n_8), .Z(n_0_704));
   MUX2_X1 i_0_0_112 (.A(\mem[8] [15]), .B(data[15]), .S(n_9), .Z(n_0_703));
   MUX2_X1 i_0_0_113 (.A(\mem[8] [14]), .B(data[14]), .S(n_9), .Z(n_0_702));
   MUX2_X1 i_0_0_114 (.A(\mem[8] [13]), .B(data[13]), .S(n_9), .Z(n_0_701));
   MUX2_X1 i_0_0_115 (.A(\mem[8] [12]), .B(data[12]), .S(n_9), .Z(n_0_700));
   MUX2_X1 i_0_0_116 (.A(\mem[8] [11]), .B(data[11]), .S(n_9), .Z(n_0_699));
   MUX2_X1 i_0_0_117 (.A(\mem[8] [10]), .B(data[10]), .S(n_9), .Z(n_0_698));
   MUX2_X1 i_0_0_118 (.A(\mem[8] [9]), .B(data[9]), .S(n_9), .Z(n_0_697));
   MUX2_X1 i_0_0_119 (.A(\mem[8] [8]), .B(data[8]), .S(n_9), .Z(n_0_696));
   MUX2_X1 i_0_0_120 (.A(\mem[8] [7]), .B(data[7]), .S(n_9), .Z(n_0_695));
   MUX2_X1 i_0_0_121 (.A(\mem[8] [6]), .B(data[6]), .S(n_9), .Z(n_0_694));
   MUX2_X1 i_0_0_122 (.A(\mem[8] [5]), .B(data[5]), .S(n_9), .Z(n_0_693));
   MUX2_X1 i_0_0_123 (.A(\mem[8] [4]), .B(data[4]), .S(n_9), .Z(n_0_692));
   MUX2_X1 i_0_0_124 (.A(\mem[8] [3]), .B(data[3]), .S(n_9), .Z(n_0_691));
   MUX2_X1 i_0_0_125 (.A(\mem[8] [2]), .B(data[2]), .S(n_9), .Z(n_0_690));
   MUX2_X1 i_0_0_126 (.A(\mem[8] [1]), .B(data[1]), .S(n_9), .Z(n_0_689));
   MUX2_X1 i_0_0_127 (.A(\mem[8] [0]), .B(data[0]), .S(n_9), .Z(n_0_688));
   MUX2_X1 i_0_0_128 (.A(\mem[9] [15]), .B(data[15]), .S(n_10), .Z(n_0_687));
   MUX2_X1 i_0_0_129 (.A(\mem[9] [14]), .B(data[14]), .S(n_10), .Z(n_0_686));
   MUX2_X1 i_0_0_130 (.A(\mem[9] [13]), .B(data[13]), .S(n_10), .Z(n_0_685));
   MUX2_X1 i_0_0_131 (.A(\mem[9] [12]), .B(data[12]), .S(n_10), .Z(n_0_684));
   MUX2_X1 i_0_0_132 (.A(\mem[9] [11]), .B(data[11]), .S(n_10), .Z(n_0_683));
   MUX2_X1 i_0_0_133 (.A(\mem[9] [10]), .B(data[10]), .S(n_10), .Z(n_0_682));
   MUX2_X1 i_0_0_134 (.A(\mem[9] [9]), .B(data[9]), .S(n_10), .Z(n_0_681));
   MUX2_X1 i_0_0_135 (.A(\mem[9] [8]), .B(data[8]), .S(n_10), .Z(n_0_680));
   MUX2_X1 i_0_0_136 (.A(\mem[9] [7]), .B(data[7]), .S(n_10), .Z(n_0_679));
   MUX2_X1 i_0_0_137 (.A(\mem[9] [6]), .B(data[6]), .S(n_10), .Z(n_0_678));
   MUX2_X1 i_0_0_138 (.A(\mem[9] [5]), .B(data[5]), .S(n_10), .Z(n_0_677));
   MUX2_X1 i_0_0_139 (.A(\mem[9] [4]), .B(data[4]), .S(n_10), .Z(n_0_676));
   MUX2_X1 i_0_0_140 (.A(\mem[9] [3]), .B(data[3]), .S(n_10), .Z(n_0_675));
   MUX2_X1 i_0_0_141 (.A(\mem[9] [2]), .B(data[2]), .S(n_10), .Z(n_0_674));
   MUX2_X1 i_0_0_142 (.A(\mem[9] [1]), .B(data[1]), .S(n_10), .Z(n_0_673));
   MUX2_X1 i_0_0_143 (.A(\mem[9] [0]), .B(data[0]), .S(n_10), .Z(n_0_672));
   MUX2_X1 i_0_0_144 (.A(\mem[10] [15]), .B(data[15]), .S(n_11), .Z(n_0_671));
   MUX2_X1 i_0_0_145 (.A(\mem[10] [14]), .B(data[14]), .S(n_11), .Z(n_0_670));
   MUX2_X1 i_0_0_146 (.A(\mem[10] [13]), .B(data[13]), .S(n_11), .Z(n_0_669));
   MUX2_X1 i_0_0_147 (.A(\mem[10] [12]), .B(data[12]), .S(n_11), .Z(n_0_668));
   MUX2_X1 i_0_0_148 (.A(\mem[10] [11]), .B(data[11]), .S(n_11), .Z(n_0_667));
   MUX2_X1 i_0_0_149 (.A(\mem[10] [10]), .B(data[10]), .S(n_11), .Z(n_0_666));
   MUX2_X1 i_0_0_150 (.A(\mem[10] [9]), .B(data[9]), .S(n_11), .Z(n_0_665));
   MUX2_X1 i_0_0_151 (.A(\mem[10] [8]), .B(data[8]), .S(n_11), .Z(n_0_664));
   MUX2_X1 i_0_0_152 (.A(\mem[10] [7]), .B(data[7]), .S(n_11), .Z(n_0_663));
   MUX2_X1 i_0_0_153 (.A(\mem[10] [6]), .B(data[6]), .S(n_11), .Z(n_0_662));
   MUX2_X1 i_0_0_154 (.A(\mem[10] [5]), .B(data[5]), .S(n_11), .Z(n_0_661));
   MUX2_X1 i_0_0_155 (.A(\mem[10] [4]), .B(data[4]), .S(n_11), .Z(n_0_660));
   MUX2_X1 i_0_0_156 (.A(\mem[10] [3]), .B(data[3]), .S(n_11), .Z(n_0_659));
   MUX2_X1 i_0_0_157 (.A(\mem[10] [2]), .B(data[2]), .S(n_11), .Z(n_0_658));
   MUX2_X1 i_0_0_158 (.A(\mem[10] [1]), .B(data[1]), .S(n_11), .Z(n_0_657));
   MUX2_X1 i_0_0_159 (.A(\mem[10] [0]), .B(data[0]), .S(n_11), .Z(n_0_656));
   MUX2_X1 i_0_0_160 (.A(\mem[11] [15]), .B(data[15]), .S(n_12), .Z(n_0_655));
   MUX2_X1 i_0_0_161 (.A(\mem[11] [14]), .B(data[14]), .S(n_12), .Z(n_0_654));
   MUX2_X1 i_0_0_162 (.A(\mem[11] [13]), .B(data[13]), .S(n_12), .Z(n_0_653));
   MUX2_X1 i_0_0_163 (.A(\mem[11] [12]), .B(data[12]), .S(n_12), .Z(n_0_652));
   MUX2_X1 i_0_0_164 (.A(\mem[11] [11]), .B(data[11]), .S(n_12), .Z(n_0_651));
   MUX2_X1 i_0_0_165 (.A(\mem[11] [10]), .B(data[10]), .S(n_12), .Z(n_0_650));
   MUX2_X1 i_0_0_166 (.A(\mem[11] [9]), .B(data[9]), .S(n_12), .Z(n_0_649));
   MUX2_X1 i_0_0_167 (.A(\mem[11] [8]), .B(data[8]), .S(n_12), .Z(n_0_648));
   MUX2_X1 i_0_0_168 (.A(\mem[11] [7]), .B(data[7]), .S(n_12), .Z(n_0_647));
   MUX2_X1 i_0_0_169 (.A(\mem[11] [6]), .B(data[6]), .S(n_12), .Z(n_0_646));
   MUX2_X1 i_0_0_170 (.A(\mem[11] [5]), .B(data[5]), .S(n_12), .Z(n_0_645));
   MUX2_X1 i_0_0_171 (.A(\mem[11] [4]), .B(data[4]), .S(n_12), .Z(n_0_644));
   MUX2_X1 i_0_0_172 (.A(\mem[11] [3]), .B(data[3]), .S(n_12), .Z(n_0_643));
   MUX2_X1 i_0_0_173 (.A(\mem[11] [2]), .B(data[2]), .S(n_12), .Z(n_0_642));
   MUX2_X1 i_0_0_174 (.A(\mem[11] [1]), .B(data[1]), .S(n_12), .Z(n_0_641));
   MUX2_X1 i_0_0_175 (.A(\mem[11] [0]), .B(data[0]), .S(n_12), .Z(n_0_640));
   MUX2_X1 i_0_0_176 (.A(\mem[12] [15]), .B(data[15]), .S(n_13), .Z(n_0_639));
   MUX2_X1 i_0_0_177 (.A(\mem[12] [14]), .B(data[14]), .S(n_13), .Z(n_0_638));
   MUX2_X1 i_0_0_178 (.A(\mem[12] [13]), .B(data[13]), .S(n_13), .Z(n_0_637));
   MUX2_X1 i_0_0_179 (.A(\mem[12] [12]), .B(data[12]), .S(n_13), .Z(n_0_636));
   MUX2_X1 i_0_0_180 (.A(\mem[12] [11]), .B(data[11]), .S(n_13), .Z(n_0_635));
   MUX2_X1 i_0_0_181 (.A(\mem[12] [10]), .B(data[10]), .S(n_13), .Z(n_0_634));
   MUX2_X1 i_0_0_182 (.A(\mem[12] [9]), .B(data[9]), .S(n_13), .Z(n_0_633));
   MUX2_X1 i_0_0_183 (.A(\mem[12] [8]), .B(data[8]), .S(n_13), .Z(n_0_632));
   MUX2_X1 i_0_0_184 (.A(\mem[12] [7]), .B(data[7]), .S(n_13), .Z(n_0_631));
   MUX2_X1 i_0_0_185 (.A(\mem[12] [6]), .B(data[6]), .S(n_13), .Z(n_0_630));
   MUX2_X1 i_0_0_186 (.A(\mem[12] [5]), .B(data[5]), .S(n_13), .Z(n_0_629));
   MUX2_X1 i_0_0_187 (.A(\mem[12] [4]), .B(data[4]), .S(n_13), .Z(n_0_628));
   MUX2_X1 i_0_0_188 (.A(\mem[12] [3]), .B(data[3]), .S(n_13), .Z(n_0_627));
   MUX2_X1 i_0_0_189 (.A(\mem[12] [2]), .B(data[2]), .S(n_13), .Z(n_0_626));
   MUX2_X1 i_0_0_190 (.A(\mem[12] [1]), .B(data[1]), .S(n_13), .Z(n_0_625));
   MUX2_X1 i_0_0_191 (.A(\mem[12] [0]), .B(data[0]), .S(n_13), .Z(n_0_624));
   MUX2_X1 i_0_0_192 (.A(\mem[13] [15]), .B(data[15]), .S(n_14), .Z(n_0_623));
   MUX2_X1 i_0_0_193 (.A(\mem[13] [14]), .B(data[14]), .S(n_14), .Z(n_0_622));
   MUX2_X1 i_0_0_194 (.A(\mem[13] [13]), .B(data[13]), .S(n_14), .Z(n_0_621));
   MUX2_X1 i_0_0_195 (.A(\mem[13] [12]), .B(data[12]), .S(n_14), .Z(n_0_620));
   MUX2_X1 i_0_0_196 (.A(\mem[13] [11]), .B(data[11]), .S(n_14), .Z(n_0_619));
   MUX2_X1 i_0_0_197 (.A(\mem[13] [10]), .B(data[10]), .S(n_14), .Z(n_0_618));
   MUX2_X1 i_0_0_198 (.A(\mem[13] [9]), .B(data[9]), .S(n_14), .Z(n_0_617));
   MUX2_X1 i_0_0_199 (.A(\mem[13] [8]), .B(data[8]), .S(n_14), .Z(n_0_616));
   MUX2_X1 i_0_0_200 (.A(\mem[13] [7]), .B(data[7]), .S(n_14), .Z(n_0_615));
   MUX2_X1 i_0_0_201 (.A(\mem[13] [6]), .B(data[6]), .S(n_14), .Z(n_0_614));
   MUX2_X1 i_0_0_202 (.A(\mem[13] [5]), .B(data[5]), .S(n_14), .Z(n_0_613));
   MUX2_X1 i_0_0_203 (.A(\mem[13] [4]), .B(data[4]), .S(n_14), .Z(n_0_612));
   MUX2_X1 i_0_0_204 (.A(\mem[13] [3]), .B(data[3]), .S(n_14), .Z(n_0_611));
   MUX2_X1 i_0_0_205 (.A(\mem[13] [2]), .B(data[2]), .S(n_14), .Z(n_0_610));
   MUX2_X1 i_0_0_206 (.A(\mem[13] [1]), .B(data[1]), .S(n_14), .Z(n_0_609));
   MUX2_X1 i_0_0_207 (.A(\mem[13] [0]), .B(data[0]), .S(n_14), .Z(n_0_608));
   MUX2_X1 i_0_0_208 (.A(\mem[14] [15]), .B(data[15]), .S(n_15), .Z(n_0_607));
   MUX2_X1 i_0_0_209 (.A(\mem[14] [14]), .B(data[14]), .S(n_15), .Z(n_0_606));
   MUX2_X1 i_0_0_210 (.A(\mem[14] [13]), .B(data[13]), .S(n_15), .Z(n_0_605));
   MUX2_X1 i_0_0_211 (.A(\mem[14] [12]), .B(data[12]), .S(n_15), .Z(n_0_604));
   MUX2_X1 i_0_0_212 (.A(\mem[14] [11]), .B(data[11]), .S(n_15), .Z(n_0_603));
   MUX2_X1 i_0_0_213 (.A(\mem[14] [10]), .B(data[10]), .S(n_15), .Z(n_0_602));
   MUX2_X1 i_0_0_214 (.A(\mem[14] [9]), .B(data[9]), .S(n_15), .Z(n_0_601));
   MUX2_X1 i_0_0_215 (.A(\mem[14] [8]), .B(data[8]), .S(n_15), .Z(n_0_600));
   MUX2_X1 i_0_0_216 (.A(\mem[14] [7]), .B(data[7]), .S(n_15), .Z(n_0_599));
   MUX2_X1 i_0_0_217 (.A(\mem[14] [6]), .B(data[6]), .S(n_15), .Z(n_0_598));
   MUX2_X1 i_0_0_218 (.A(\mem[14] [5]), .B(data[5]), .S(n_15), .Z(n_0_597));
   MUX2_X1 i_0_0_219 (.A(\mem[14] [4]), .B(data[4]), .S(n_15), .Z(n_0_596));
   MUX2_X1 i_0_0_220 (.A(\mem[14] [3]), .B(data[3]), .S(n_15), .Z(n_0_595));
   MUX2_X1 i_0_0_221 (.A(\mem[14] [2]), .B(data[2]), .S(n_15), .Z(n_0_594));
   MUX2_X1 i_0_0_222 (.A(\mem[14] [1]), .B(data[1]), .S(n_15), .Z(n_0_593));
   MUX2_X1 i_0_0_223 (.A(\mem[14] [0]), .B(data[0]), .S(n_15), .Z(n_0_592));
   MUX2_X1 i_0_0_224 (.A(\mem[15] [15]), .B(data[15]), .S(n_16), .Z(n_0_591));
   MUX2_X1 i_0_0_225 (.A(\mem[15] [14]), .B(data[14]), .S(n_16), .Z(n_0_590));
   MUX2_X1 i_0_0_226 (.A(\mem[15] [13]), .B(data[13]), .S(n_16), .Z(n_0_589));
   MUX2_X1 i_0_0_227 (.A(\mem[15] [12]), .B(data[12]), .S(n_16), .Z(n_0_588));
   MUX2_X1 i_0_0_228 (.A(\mem[15] [11]), .B(data[11]), .S(n_16), .Z(n_0_587));
   MUX2_X1 i_0_0_229 (.A(\mem[15] [10]), .B(data[10]), .S(n_16), .Z(n_0_586));
   MUX2_X1 i_0_0_230 (.A(\mem[15] [9]), .B(data[9]), .S(n_16), .Z(n_0_585));
   MUX2_X1 i_0_0_231 (.A(\mem[15] [8]), .B(data[8]), .S(n_16), .Z(n_0_584));
   MUX2_X1 i_0_0_232 (.A(\mem[15] [7]), .B(data[7]), .S(n_16), .Z(n_0_583));
   MUX2_X1 i_0_0_233 (.A(\mem[15] [6]), .B(data[6]), .S(n_16), .Z(n_0_582));
   MUX2_X1 i_0_0_234 (.A(\mem[15] [5]), .B(data[5]), .S(n_16), .Z(n_0_581));
   MUX2_X1 i_0_0_235 (.A(\mem[15] [4]), .B(data[4]), .S(n_16), .Z(n_0_580));
   MUX2_X1 i_0_0_236 (.A(\mem[15] [3]), .B(data[3]), .S(n_16), .Z(n_0_579));
   MUX2_X1 i_0_0_237 (.A(\mem[15] [2]), .B(data[2]), .S(n_16), .Z(n_0_578));
   MUX2_X1 i_0_0_238 (.A(\mem[15] [1]), .B(data[1]), .S(n_16), .Z(n_0_577));
   MUX2_X1 i_0_0_239 (.A(\mem[15] [0]), .B(data[0]), .S(n_16), .Z(n_0_576));
   MUX2_X1 i_0_0_240 (.A(\mem[16] [15]), .B(data[15]), .S(n_17), .Z(n_0_575));
   MUX2_X1 i_0_0_241 (.A(\mem[16] [14]), .B(data[14]), .S(n_17), .Z(n_0_574));
   MUX2_X1 i_0_0_242 (.A(\mem[16] [13]), .B(data[13]), .S(n_17), .Z(n_0_573));
   MUX2_X1 i_0_0_243 (.A(\mem[16] [12]), .B(data[12]), .S(n_17), .Z(n_0_572));
   MUX2_X1 i_0_0_244 (.A(\mem[16] [11]), .B(data[11]), .S(n_17), .Z(n_0_571));
   MUX2_X1 i_0_0_245 (.A(\mem[16] [10]), .B(data[10]), .S(n_17), .Z(n_0_570));
   MUX2_X1 i_0_0_246 (.A(\mem[16] [9]), .B(data[9]), .S(n_17), .Z(n_0_569));
   MUX2_X1 i_0_0_247 (.A(\mem[16] [8]), .B(data[8]), .S(n_17), .Z(n_0_568));
   MUX2_X1 i_0_0_248 (.A(\mem[16] [7]), .B(data[7]), .S(n_17), .Z(n_0_567));
   MUX2_X1 i_0_0_249 (.A(\mem[16] [6]), .B(data[6]), .S(n_17), .Z(n_0_566));
   MUX2_X1 i_0_0_250 (.A(\mem[16] [5]), .B(data[5]), .S(n_17), .Z(n_0_565));
   MUX2_X1 i_0_0_251 (.A(\mem[16] [4]), .B(data[4]), .S(n_17), .Z(n_0_564));
   MUX2_X1 i_0_0_252 (.A(\mem[16] [3]), .B(data[3]), .S(n_17), .Z(n_0_563));
   MUX2_X1 i_0_0_253 (.A(\mem[16] [2]), .B(data[2]), .S(n_17), .Z(n_0_562));
   MUX2_X1 i_0_0_254 (.A(\mem[16] [1]), .B(data[1]), .S(n_17), .Z(n_0_561));
   MUX2_X1 i_0_0_255 (.A(\mem[16] [0]), .B(data[0]), .S(n_17), .Z(n_0_560));
   MUX2_X1 i_0_0_256 (.A(\mem[17] [15]), .B(data[15]), .S(n_18), .Z(n_0_559));
   MUX2_X1 i_0_0_257 (.A(\mem[17] [14]), .B(data[14]), .S(n_18), .Z(n_0_558));
   MUX2_X1 i_0_0_258 (.A(\mem[17] [13]), .B(data[13]), .S(n_18), .Z(n_0_557));
   MUX2_X1 i_0_0_259 (.A(\mem[17] [12]), .B(data[12]), .S(n_18), .Z(n_0_556));
   MUX2_X1 i_0_0_260 (.A(\mem[17] [11]), .B(data[11]), .S(n_18), .Z(n_0_555));
   MUX2_X1 i_0_0_261 (.A(\mem[17] [10]), .B(data[10]), .S(n_18), .Z(n_0_554));
   MUX2_X1 i_0_0_262 (.A(\mem[17] [9]), .B(data[9]), .S(n_18), .Z(n_0_553));
   MUX2_X1 i_0_0_263 (.A(\mem[17] [8]), .B(data[8]), .S(n_18), .Z(n_0_552));
   MUX2_X1 i_0_0_264 (.A(\mem[17] [7]), .B(data[7]), .S(n_18), .Z(n_0_551));
   MUX2_X1 i_0_0_265 (.A(\mem[17] [6]), .B(data[6]), .S(n_18), .Z(n_0_550));
   MUX2_X1 i_0_0_266 (.A(\mem[17] [5]), .B(data[5]), .S(n_18), .Z(n_0_549));
   MUX2_X1 i_0_0_267 (.A(\mem[17] [4]), .B(data[4]), .S(n_18), .Z(n_0_548));
   MUX2_X1 i_0_0_268 (.A(\mem[17] [3]), .B(data[3]), .S(n_18), .Z(n_0_547));
   MUX2_X1 i_0_0_269 (.A(\mem[17] [2]), .B(data[2]), .S(n_18), .Z(n_0_546));
   MUX2_X1 i_0_0_270 (.A(\mem[17] [1]), .B(data[1]), .S(n_18), .Z(n_0_545));
   MUX2_X1 i_0_0_271 (.A(\mem[17] [0]), .B(data[0]), .S(n_18), .Z(n_0_544));
   MUX2_X1 i_0_0_272 (.A(\mem[18] [15]), .B(data[15]), .S(n_19), .Z(n_0_543));
   MUX2_X1 i_0_0_273 (.A(\mem[18] [14]), .B(data[14]), .S(n_19), .Z(n_0_542));
   MUX2_X1 i_0_0_274 (.A(\mem[18] [13]), .B(data[13]), .S(n_19), .Z(n_0_541));
   MUX2_X1 i_0_0_275 (.A(\mem[18] [12]), .B(data[12]), .S(n_19), .Z(n_0_540));
   MUX2_X1 i_0_0_276 (.A(\mem[18] [11]), .B(data[11]), .S(n_19), .Z(n_0_539));
   MUX2_X1 i_0_0_277 (.A(\mem[18] [10]), .B(data[10]), .S(n_19), .Z(n_0_538));
   MUX2_X1 i_0_0_278 (.A(\mem[18] [9]), .B(data[9]), .S(n_19), .Z(n_0_537));
   MUX2_X1 i_0_0_279 (.A(\mem[18] [8]), .B(data[8]), .S(n_19), .Z(n_0_536));
   MUX2_X1 i_0_0_280 (.A(\mem[18] [7]), .B(data[7]), .S(n_19), .Z(n_0_535));
   MUX2_X1 i_0_0_281 (.A(\mem[18] [6]), .B(data[6]), .S(n_19), .Z(n_0_534));
   MUX2_X1 i_0_0_282 (.A(\mem[18] [5]), .B(data[5]), .S(n_19), .Z(n_0_533));
   MUX2_X1 i_0_0_283 (.A(\mem[18] [4]), .B(data[4]), .S(n_19), .Z(n_0_532));
   MUX2_X1 i_0_0_284 (.A(\mem[18] [3]), .B(data[3]), .S(n_19), .Z(n_0_531));
   MUX2_X1 i_0_0_285 (.A(\mem[18] [2]), .B(data[2]), .S(n_19), .Z(n_0_530));
   MUX2_X1 i_0_0_286 (.A(\mem[18] [1]), .B(data[1]), .S(n_19), .Z(n_0_529));
   MUX2_X1 i_0_0_287 (.A(\mem[18] [0]), .B(data[0]), .S(n_19), .Z(n_0_528));
   MUX2_X1 i_0_0_288 (.A(\mem[19] [15]), .B(data[15]), .S(n_20), .Z(n_0_527));
   MUX2_X1 i_0_0_289 (.A(\mem[19] [14]), .B(data[14]), .S(n_20), .Z(n_0_526));
   MUX2_X1 i_0_0_290 (.A(\mem[19] [13]), .B(data[13]), .S(n_20), .Z(n_0_525));
   MUX2_X1 i_0_0_291 (.A(\mem[19] [12]), .B(data[12]), .S(n_20), .Z(n_0_524));
   MUX2_X1 i_0_0_292 (.A(\mem[19] [11]), .B(data[11]), .S(n_20), .Z(n_0_523));
   MUX2_X1 i_0_0_293 (.A(\mem[19] [10]), .B(data[10]), .S(n_20), .Z(n_0_522));
   MUX2_X1 i_0_0_294 (.A(\mem[19] [9]), .B(data[9]), .S(n_20), .Z(n_0_521));
   MUX2_X1 i_0_0_295 (.A(\mem[19] [8]), .B(data[8]), .S(n_20), .Z(n_0_520));
   MUX2_X1 i_0_0_296 (.A(\mem[19] [7]), .B(data[7]), .S(n_20), .Z(n_0_519));
   MUX2_X1 i_0_0_297 (.A(\mem[19] [6]), .B(data[6]), .S(n_20), .Z(n_0_518));
   MUX2_X1 i_0_0_298 (.A(\mem[19] [5]), .B(data[5]), .S(n_20), .Z(n_0_517));
   MUX2_X1 i_0_0_299 (.A(\mem[19] [4]), .B(data[4]), .S(n_20), .Z(n_0_516));
   MUX2_X1 i_0_0_300 (.A(\mem[19] [3]), .B(data[3]), .S(n_20), .Z(n_0_515));
   MUX2_X1 i_0_0_301 (.A(\mem[19] [2]), .B(data[2]), .S(n_20), .Z(n_0_514));
   MUX2_X1 i_0_0_302 (.A(\mem[19] [1]), .B(data[1]), .S(n_20), .Z(n_0_513));
   MUX2_X1 i_0_0_303 (.A(\mem[19] [0]), .B(data[0]), .S(n_20), .Z(n_0_512));
   MUX2_X1 i_0_0_304 (.A(\mem[20] [15]), .B(data[15]), .S(n_21), .Z(n_0_511));
   MUX2_X1 i_0_0_305 (.A(\mem[20] [14]), .B(data[14]), .S(n_21), .Z(n_0_510));
   MUX2_X1 i_0_0_306 (.A(\mem[20] [13]), .B(data[13]), .S(n_21), .Z(n_0_509));
   MUX2_X1 i_0_0_307 (.A(\mem[20] [12]), .B(data[12]), .S(n_21), .Z(n_0_508));
   MUX2_X1 i_0_0_308 (.A(\mem[20] [11]), .B(data[11]), .S(n_21), .Z(n_0_507));
   MUX2_X1 i_0_0_309 (.A(\mem[20] [10]), .B(data[10]), .S(n_21), .Z(n_0_506));
   MUX2_X1 i_0_0_310 (.A(\mem[20] [9]), .B(data[9]), .S(n_21), .Z(n_0_505));
   MUX2_X1 i_0_0_311 (.A(\mem[20] [8]), .B(data[8]), .S(n_21), .Z(n_0_504));
   MUX2_X1 i_0_0_312 (.A(\mem[20] [7]), .B(data[7]), .S(n_21), .Z(n_0_503));
   MUX2_X1 i_0_0_313 (.A(\mem[20] [6]), .B(data[6]), .S(n_21), .Z(n_0_502));
   MUX2_X1 i_0_0_314 (.A(\mem[20] [5]), .B(data[5]), .S(n_21), .Z(n_0_501));
   MUX2_X1 i_0_0_315 (.A(\mem[20] [4]), .B(data[4]), .S(n_21), .Z(n_0_500));
   MUX2_X1 i_0_0_316 (.A(\mem[20] [3]), .B(data[3]), .S(n_21), .Z(n_0_499));
   MUX2_X1 i_0_0_317 (.A(\mem[20] [2]), .B(data[2]), .S(n_21), .Z(n_0_498));
   MUX2_X1 i_0_0_318 (.A(\mem[20] [1]), .B(data[1]), .S(n_21), .Z(n_0_497));
   MUX2_X1 i_0_0_319 (.A(\mem[20] [0]), .B(data[0]), .S(n_21), .Z(n_0_496));
   MUX2_X1 i_0_0_320 (.A(\mem[21] [15]), .B(data[15]), .S(n_22), .Z(n_0_495));
   MUX2_X1 i_0_0_321 (.A(\mem[21] [14]), .B(data[14]), .S(n_22), .Z(n_0_494));
   MUX2_X1 i_0_0_322 (.A(\mem[21] [13]), .B(data[13]), .S(n_22), .Z(n_0_493));
   MUX2_X1 i_0_0_323 (.A(\mem[21] [12]), .B(data[12]), .S(n_22), .Z(n_0_492));
   MUX2_X1 i_0_0_324 (.A(\mem[21] [11]), .B(data[11]), .S(n_22), .Z(n_0_491));
   MUX2_X1 i_0_0_325 (.A(\mem[21] [10]), .B(data[10]), .S(n_22), .Z(n_0_490));
   MUX2_X1 i_0_0_326 (.A(\mem[21] [9]), .B(data[9]), .S(n_22), .Z(n_0_489));
   MUX2_X1 i_0_0_327 (.A(\mem[21] [8]), .B(data[8]), .S(n_22), .Z(n_0_488));
   MUX2_X1 i_0_0_328 (.A(\mem[21] [7]), .B(data[7]), .S(n_22), .Z(n_0_487));
   MUX2_X1 i_0_0_329 (.A(\mem[21] [6]), .B(data[6]), .S(n_22), .Z(n_0_486));
   MUX2_X1 i_0_0_330 (.A(\mem[21] [5]), .B(data[5]), .S(n_22), .Z(n_0_485));
   MUX2_X1 i_0_0_331 (.A(\mem[21] [4]), .B(data[4]), .S(n_22), .Z(n_0_484));
   MUX2_X1 i_0_0_332 (.A(\mem[21] [3]), .B(data[3]), .S(n_22), .Z(n_0_483));
   MUX2_X1 i_0_0_333 (.A(\mem[21] [2]), .B(data[2]), .S(n_22), .Z(n_0_482));
   MUX2_X1 i_0_0_334 (.A(\mem[21] [1]), .B(data[1]), .S(n_22), .Z(n_0_481));
   MUX2_X1 i_0_0_335 (.A(\mem[21] [0]), .B(data[0]), .S(n_22), .Z(n_0_480));
   MUX2_X1 i_0_0_336 (.A(\mem[22] [15]), .B(data[15]), .S(n_23), .Z(n_0_479));
   MUX2_X1 i_0_0_337 (.A(\mem[22] [14]), .B(data[14]), .S(n_23), .Z(n_0_478));
   MUX2_X1 i_0_0_338 (.A(\mem[22] [13]), .B(data[13]), .S(n_23), .Z(n_0_477));
   MUX2_X1 i_0_0_339 (.A(\mem[22] [12]), .B(data[12]), .S(n_23), .Z(n_0_476));
   MUX2_X1 i_0_0_340 (.A(\mem[22] [11]), .B(data[11]), .S(n_23), .Z(n_0_475));
   MUX2_X1 i_0_0_341 (.A(\mem[22] [10]), .B(data[10]), .S(n_23), .Z(n_0_474));
   MUX2_X1 i_0_0_342 (.A(\mem[22] [9]), .B(data[9]), .S(n_23), .Z(n_0_473));
   MUX2_X1 i_0_0_343 (.A(\mem[22] [8]), .B(data[8]), .S(n_23), .Z(n_0_472));
   MUX2_X1 i_0_0_344 (.A(\mem[22] [7]), .B(data[7]), .S(n_23), .Z(n_0_471));
   MUX2_X1 i_0_0_345 (.A(\mem[22] [6]), .B(data[6]), .S(n_23), .Z(n_0_470));
   MUX2_X1 i_0_0_346 (.A(\mem[22] [5]), .B(data[5]), .S(n_23), .Z(n_0_469));
   MUX2_X1 i_0_0_347 (.A(\mem[22] [4]), .B(data[4]), .S(n_23), .Z(n_0_468));
   MUX2_X1 i_0_0_348 (.A(\mem[22] [3]), .B(data[3]), .S(n_23), .Z(n_0_467));
   MUX2_X1 i_0_0_349 (.A(\mem[22] [2]), .B(data[2]), .S(n_23), .Z(n_0_466));
   MUX2_X1 i_0_0_350 (.A(\mem[22] [1]), .B(data[1]), .S(n_23), .Z(n_0_465));
   MUX2_X1 i_0_0_351 (.A(\mem[22] [0]), .B(data[0]), .S(n_23), .Z(n_0_464));
   MUX2_X1 i_0_0_352 (.A(\mem[23] [15]), .B(data[15]), .S(n_24), .Z(n_0_463));
   MUX2_X1 i_0_0_353 (.A(\mem[23] [14]), .B(data[14]), .S(n_24), .Z(n_0_462));
   MUX2_X1 i_0_0_354 (.A(\mem[23] [13]), .B(data[13]), .S(n_24), .Z(n_0_461));
   MUX2_X1 i_0_0_355 (.A(\mem[23] [12]), .B(data[12]), .S(n_24), .Z(n_0_460));
   MUX2_X1 i_0_0_356 (.A(\mem[23] [11]), .B(data[11]), .S(n_24), .Z(n_0_459));
   MUX2_X1 i_0_0_357 (.A(\mem[23] [10]), .B(data[10]), .S(n_24), .Z(n_0_458));
   MUX2_X1 i_0_0_358 (.A(\mem[23] [9]), .B(data[9]), .S(n_24), .Z(n_0_457));
   MUX2_X1 i_0_0_359 (.A(\mem[23] [8]), .B(data[8]), .S(n_24), .Z(n_0_456));
   MUX2_X1 i_0_0_360 (.A(\mem[23] [7]), .B(data[7]), .S(n_24), .Z(n_0_455));
   MUX2_X1 i_0_0_361 (.A(\mem[23] [6]), .B(data[6]), .S(n_24), .Z(n_0_454));
   MUX2_X1 i_0_0_362 (.A(\mem[23] [5]), .B(data[5]), .S(n_24), .Z(n_0_453));
   MUX2_X1 i_0_0_363 (.A(\mem[23] [4]), .B(data[4]), .S(n_24), .Z(n_0_452));
   MUX2_X1 i_0_0_364 (.A(\mem[23] [3]), .B(data[3]), .S(n_24), .Z(n_0_451));
   MUX2_X1 i_0_0_365 (.A(\mem[23] [2]), .B(data[2]), .S(n_24), .Z(n_0_450));
   MUX2_X1 i_0_0_366 (.A(\mem[23] [1]), .B(data[1]), .S(n_24), .Z(n_0_449));
   MUX2_X1 i_0_0_367 (.A(\mem[23] [0]), .B(data[0]), .S(n_24), .Z(n_0_448));
   MUX2_X1 i_0_0_368 (.A(\mem[24] [15]), .B(data[15]), .S(n_25), .Z(n_0_447));
   MUX2_X1 i_0_0_369 (.A(\mem[24] [14]), .B(data[14]), .S(n_25), .Z(n_0_446));
   MUX2_X1 i_0_0_370 (.A(\mem[24] [13]), .B(data[13]), .S(n_25), .Z(n_0_445));
   MUX2_X1 i_0_0_371 (.A(\mem[24] [12]), .B(data[12]), .S(n_25), .Z(n_0_444));
   MUX2_X1 i_0_0_372 (.A(\mem[24] [11]), .B(data[11]), .S(n_25), .Z(n_0_443));
   MUX2_X1 i_0_0_373 (.A(\mem[24] [10]), .B(data[10]), .S(n_25), .Z(n_0_442));
   MUX2_X1 i_0_0_374 (.A(\mem[24] [9]), .B(data[9]), .S(n_25), .Z(n_0_441));
   MUX2_X1 i_0_0_375 (.A(\mem[24] [8]), .B(data[8]), .S(n_25), .Z(n_0_440));
   MUX2_X1 i_0_0_376 (.A(\mem[24] [7]), .B(data[7]), .S(n_25), .Z(n_0_439));
   MUX2_X1 i_0_0_377 (.A(\mem[24] [6]), .B(data[6]), .S(n_25), .Z(n_0_438));
   MUX2_X1 i_0_0_378 (.A(\mem[24] [5]), .B(data[5]), .S(n_25), .Z(n_0_437));
   MUX2_X1 i_0_0_379 (.A(\mem[24] [4]), .B(data[4]), .S(n_25), .Z(n_0_436));
   MUX2_X1 i_0_0_380 (.A(\mem[24] [3]), .B(data[3]), .S(n_25), .Z(n_0_435));
   MUX2_X1 i_0_0_381 (.A(\mem[24] [2]), .B(data[2]), .S(n_25), .Z(n_0_434));
   MUX2_X1 i_0_0_382 (.A(\mem[24] [1]), .B(data[1]), .S(n_25), .Z(n_0_433));
   MUX2_X1 i_0_0_383 (.A(\mem[24] [0]), .B(data[0]), .S(n_25), .Z(n_0_432));
   MUX2_X1 i_0_0_384 (.A(\mem[25] [15]), .B(data[15]), .S(n_26), .Z(n_0_431));
   MUX2_X1 i_0_0_385 (.A(\mem[25] [14]), .B(data[14]), .S(n_26), .Z(n_0_430));
   MUX2_X1 i_0_0_386 (.A(\mem[25] [13]), .B(data[13]), .S(n_26), .Z(n_0_429));
   MUX2_X1 i_0_0_387 (.A(\mem[25] [12]), .B(data[12]), .S(n_26), .Z(n_0_428));
   MUX2_X1 i_0_0_388 (.A(\mem[25] [11]), .B(data[11]), .S(n_26), .Z(n_0_427));
   MUX2_X1 i_0_0_389 (.A(\mem[25] [10]), .B(data[10]), .S(n_26), .Z(n_0_426));
   MUX2_X1 i_0_0_390 (.A(\mem[25] [9]), .B(data[9]), .S(n_26), .Z(n_0_425));
   MUX2_X1 i_0_0_391 (.A(\mem[25] [8]), .B(data[8]), .S(n_26), .Z(n_0_424));
   MUX2_X1 i_0_0_392 (.A(\mem[25] [7]), .B(data[7]), .S(n_26), .Z(n_0_423));
   MUX2_X1 i_0_0_393 (.A(\mem[25] [6]), .B(data[6]), .S(n_26), .Z(n_0_422));
   MUX2_X1 i_0_0_394 (.A(\mem[25] [5]), .B(data[5]), .S(n_26), .Z(n_0_421));
   MUX2_X1 i_0_0_395 (.A(\mem[25] [4]), .B(data[4]), .S(n_26), .Z(n_0_420));
   MUX2_X1 i_0_0_396 (.A(\mem[25] [3]), .B(data[3]), .S(n_26), .Z(n_0_419));
   MUX2_X1 i_0_0_397 (.A(\mem[25] [2]), .B(data[2]), .S(n_26), .Z(n_0_418));
   MUX2_X1 i_0_0_398 (.A(\mem[25] [1]), .B(data[1]), .S(n_26), .Z(n_0_417));
   MUX2_X1 i_0_0_399 (.A(\mem[25] [0]), .B(data[0]), .S(n_26), .Z(n_0_416));
   MUX2_X1 i_0_0_400 (.A(\mem[26] [15]), .B(data[15]), .S(n_27), .Z(n_0_415));
   MUX2_X1 i_0_0_401 (.A(\mem[26] [14]), .B(data[14]), .S(n_27), .Z(n_0_414));
   MUX2_X1 i_0_0_402 (.A(\mem[26] [13]), .B(data[13]), .S(n_27), .Z(n_0_413));
   MUX2_X1 i_0_0_403 (.A(\mem[26] [12]), .B(data[12]), .S(n_27), .Z(n_0_412));
   MUX2_X1 i_0_0_404 (.A(\mem[26] [11]), .B(data[11]), .S(n_27), .Z(n_0_411));
   MUX2_X1 i_0_0_405 (.A(\mem[26] [10]), .B(data[10]), .S(n_27), .Z(n_0_410));
   MUX2_X1 i_0_0_406 (.A(\mem[26] [9]), .B(data[9]), .S(n_27), .Z(n_0_409));
   MUX2_X1 i_0_0_407 (.A(\mem[26] [8]), .B(data[8]), .S(n_27), .Z(n_0_408));
   MUX2_X1 i_0_0_408 (.A(\mem[26] [7]), .B(data[7]), .S(n_27), .Z(n_0_407));
   MUX2_X1 i_0_0_409 (.A(\mem[26] [6]), .B(data[6]), .S(n_27), .Z(n_0_406));
   MUX2_X1 i_0_0_410 (.A(\mem[26] [5]), .B(data[5]), .S(n_27), .Z(n_0_405));
   MUX2_X1 i_0_0_411 (.A(\mem[26] [4]), .B(data[4]), .S(n_27), .Z(n_0_404));
   MUX2_X1 i_0_0_412 (.A(\mem[26] [3]), .B(data[3]), .S(n_27), .Z(n_0_403));
   MUX2_X1 i_0_0_413 (.A(\mem[26] [2]), .B(data[2]), .S(n_27), .Z(n_0_402));
   MUX2_X1 i_0_0_414 (.A(\mem[26] [1]), .B(data[1]), .S(n_27), .Z(n_0_401));
   MUX2_X1 i_0_0_415 (.A(\mem[26] [0]), .B(data[0]), .S(n_27), .Z(n_0_400));
   MUX2_X1 i_0_0_416 (.A(\mem[27] [15]), .B(data[15]), .S(n_28), .Z(n_0_399));
   MUX2_X1 i_0_0_417 (.A(\mem[27] [14]), .B(data[14]), .S(n_28), .Z(n_0_398));
   MUX2_X1 i_0_0_418 (.A(\mem[27] [13]), .B(data[13]), .S(n_28), .Z(n_0_397));
   MUX2_X1 i_0_0_419 (.A(\mem[27] [12]), .B(data[12]), .S(n_28), .Z(n_0_396));
   MUX2_X1 i_0_0_420 (.A(\mem[27] [11]), .B(data[11]), .S(n_28), .Z(n_0_395));
   MUX2_X1 i_0_0_421 (.A(\mem[27] [10]), .B(data[10]), .S(n_28), .Z(n_0_394));
   MUX2_X1 i_0_0_422 (.A(\mem[27] [9]), .B(data[9]), .S(n_28), .Z(n_0_393));
   MUX2_X1 i_0_0_423 (.A(\mem[27] [8]), .B(data[8]), .S(n_28), .Z(n_0_392));
   MUX2_X1 i_0_0_424 (.A(\mem[27] [7]), .B(data[7]), .S(n_28), .Z(n_0_391));
   MUX2_X1 i_0_0_425 (.A(\mem[27] [6]), .B(data[6]), .S(n_28), .Z(n_0_390));
   MUX2_X1 i_0_0_426 (.A(\mem[27] [5]), .B(data[5]), .S(n_28), .Z(n_0_389));
   MUX2_X1 i_0_0_427 (.A(\mem[27] [4]), .B(data[4]), .S(n_28), .Z(n_0_388));
   MUX2_X1 i_0_0_428 (.A(\mem[27] [3]), .B(data[3]), .S(n_28), .Z(n_0_387));
   MUX2_X1 i_0_0_429 (.A(\mem[27] [2]), .B(data[2]), .S(n_28), .Z(n_0_386));
   MUX2_X1 i_0_0_430 (.A(\mem[27] [1]), .B(data[1]), .S(n_28), .Z(n_0_385));
   MUX2_X1 i_0_0_431 (.A(\mem[27] [0]), .B(data[0]), .S(n_28), .Z(n_0_384));
   MUX2_X1 i_0_0_432 (.A(\mem[28] [15]), .B(data[15]), .S(n_29), .Z(n_0_383));
   MUX2_X1 i_0_0_433 (.A(\mem[28] [14]), .B(data[14]), .S(n_29), .Z(n_0_382));
   MUX2_X1 i_0_0_434 (.A(\mem[28] [13]), .B(data[13]), .S(n_29), .Z(n_0_381));
   MUX2_X1 i_0_0_435 (.A(\mem[28] [12]), .B(data[12]), .S(n_29), .Z(n_0_380));
   MUX2_X1 i_0_0_436 (.A(\mem[28] [11]), .B(data[11]), .S(n_29), .Z(n_0_379));
   MUX2_X1 i_0_0_437 (.A(\mem[28] [10]), .B(data[10]), .S(n_29), .Z(n_0_378));
   MUX2_X1 i_0_0_438 (.A(\mem[28] [9]), .B(data[9]), .S(n_29), .Z(n_0_377));
   MUX2_X1 i_0_0_439 (.A(\mem[28] [8]), .B(data[8]), .S(n_29), .Z(n_0_376));
   MUX2_X1 i_0_0_440 (.A(\mem[28] [7]), .B(data[7]), .S(n_29), .Z(n_0_375));
   MUX2_X1 i_0_0_441 (.A(\mem[28] [6]), .B(data[6]), .S(n_29), .Z(n_0_374));
   MUX2_X1 i_0_0_442 (.A(\mem[28] [5]), .B(data[5]), .S(n_29), .Z(n_0_373));
   MUX2_X1 i_0_0_443 (.A(\mem[28] [4]), .B(data[4]), .S(n_29), .Z(n_0_372));
   MUX2_X1 i_0_0_444 (.A(\mem[28] [3]), .B(data[3]), .S(n_29), .Z(n_0_371));
   MUX2_X1 i_0_0_445 (.A(\mem[28] [2]), .B(data[2]), .S(n_29), .Z(n_0_370));
   MUX2_X1 i_0_0_446 (.A(\mem[28] [1]), .B(data[1]), .S(n_29), .Z(n_0_369));
   MUX2_X1 i_0_0_447 (.A(\mem[28] [0]), .B(data[0]), .S(n_29), .Z(n_0_368));
   MUX2_X1 i_0_0_448 (.A(\mem[29] [15]), .B(data[15]), .S(n_30), .Z(n_0_367));
   MUX2_X1 i_0_0_449 (.A(\mem[29] [14]), .B(data[14]), .S(n_30), .Z(n_0_366));
   MUX2_X1 i_0_0_450 (.A(\mem[29] [13]), .B(data[13]), .S(n_30), .Z(n_0_365));
   MUX2_X1 i_0_0_451 (.A(\mem[29] [12]), .B(data[12]), .S(n_30), .Z(n_0_364));
   MUX2_X1 i_0_0_452 (.A(\mem[29] [11]), .B(data[11]), .S(n_30), .Z(n_0_363));
   MUX2_X1 i_0_0_453 (.A(\mem[29] [10]), .B(data[10]), .S(n_30), .Z(n_0_362));
   MUX2_X1 i_0_0_454 (.A(\mem[29] [9]), .B(data[9]), .S(n_30), .Z(n_0_361));
   MUX2_X1 i_0_0_455 (.A(\mem[29] [8]), .B(data[8]), .S(n_30), .Z(n_0_360));
   MUX2_X1 i_0_0_456 (.A(\mem[29] [7]), .B(data[7]), .S(n_30), .Z(n_0_359));
   MUX2_X1 i_0_0_457 (.A(\mem[29] [6]), .B(data[6]), .S(n_30), .Z(n_0_358));
   MUX2_X1 i_0_0_458 (.A(\mem[29] [5]), .B(data[5]), .S(n_30), .Z(n_0_357));
   MUX2_X1 i_0_0_459 (.A(\mem[29] [4]), .B(data[4]), .S(n_30), .Z(n_0_356));
   MUX2_X1 i_0_0_460 (.A(\mem[29] [3]), .B(data[3]), .S(n_30), .Z(n_0_355));
   MUX2_X1 i_0_0_461 (.A(\mem[29] [2]), .B(data[2]), .S(n_30), .Z(n_0_354));
   MUX2_X1 i_0_0_462 (.A(\mem[29] [1]), .B(data[1]), .S(n_30), .Z(n_0_353));
   MUX2_X1 i_0_0_463 (.A(\mem[29] [0]), .B(data[0]), .S(n_30), .Z(n_0_352));
   MUX2_X1 i_0_0_464 (.A(\mem[30] [15]), .B(data[15]), .S(n_31), .Z(n_0_351));
   MUX2_X1 i_0_0_465 (.A(\mem[30] [14]), .B(data[14]), .S(n_31), .Z(n_0_350));
   MUX2_X1 i_0_0_466 (.A(\mem[30] [13]), .B(data[13]), .S(n_31), .Z(n_0_349));
   MUX2_X1 i_0_0_467 (.A(\mem[30] [12]), .B(data[12]), .S(n_31), .Z(n_0_348));
   MUX2_X1 i_0_0_468 (.A(\mem[30] [11]), .B(data[11]), .S(n_31), .Z(n_0_347));
   MUX2_X1 i_0_0_469 (.A(\mem[30] [10]), .B(data[10]), .S(n_31), .Z(n_0_346));
   MUX2_X1 i_0_0_470 (.A(\mem[30] [9]), .B(data[9]), .S(n_31), .Z(n_0_345));
   MUX2_X1 i_0_0_471 (.A(\mem[30] [8]), .B(data[8]), .S(n_31), .Z(n_0_344));
   MUX2_X1 i_0_0_472 (.A(\mem[30] [7]), .B(data[7]), .S(n_31), .Z(n_0_343));
   MUX2_X1 i_0_0_473 (.A(\mem[30] [6]), .B(data[6]), .S(n_31), .Z(n_0_342));
   MUX2_X1 i_0_0_474 (.A(\mem[30] [5]), .B(data[5]), .S(n_31), .Z(n_0_341));
   MUX2_X1 i_0_0_475 (.A(\mem[30] [4]), .B(data[4]), .S(n_31), .Z(n_0_340));
   MUX2_X1 i_0_0_476 (.A(\mem[30] [3]), .B(data[3]), .S(n_31), .Z(n_0_339));
   MUX2_X1 i_0_0_477 (.A(\mem[30] [2]), .B(data[2]), .S(n_31), .Z(n_0_338));
   MUX2_X1 i_0_0_478 (.A(\mem[30] [1]), .B(data[1]), .S(n_31), .Z(n_0_337));
   MUX2_X1 i_0_0_479 (.A(\mem[30] [0]), .B(data[0]), .S(n_31), .Z(n_0_336));
   MUX2_X1 i_0_0_480 (.A(\mem[31] [15]), .B(data[15]), .S(n_32), .Z(n_0_335));
   MUX2_X1 i_0_0_481 (.A(\mem[31] [14]), .B(data[14]), .S(n_32), .Z(n_0_334));
   MUX2_X1 i_0_0_482 (.A(\mem[31] [13]), .B(data[13]), .S(n_32), .Z(n_0_333));
   MUX2_X1 i_0_0_483 (.A(\mem[31] [12]), .B(data[12]), .S(n_32), .Z(n_0_332));
   MUX2_X1 i_0_0_484 (.A(\mem[31] [11]), .B(data[11]), .S(n_32), .Z(n_0_331));
   MUX2_X1 i_0_0_485 (.A(\mem[31] [10]), .B(data[10]), .S(n_32), .Z(n_0_330));
   MUX2_X1 i_0_0_486 (.A(\mem[31] [9]), .B(data[9]), .S(n_32), .Z(n_0_329));
   MUX2_X1 i_0_0_487 (.A(\mem[31] [8]), .B(data[8]), .S(n_32), .Z(n_0_328));
   MUX2_X1 i_0_0_488 (.A(\mem[31] [7]), .B(data[7]), .S(n_32), .Z(n_0_327));
   MUX2_X1 i_0_0_489 (.A(\mem[31] [6]), .B(data[6]), .S(n_32), .Z(n_0_326));
   MUX2_X1 i_0_0_490 (.A(\mem[31] [5]), .B(data[5]), .S(n_32), .Z(n_0_325));
   MUX2_X1 i_0_0_491 (.A(\mem[31] [4]), .B(data[4]), .S(n_32), .Z(n_0_324));
   MUX2_X1 i_0_0_492 (.A(\mem[31] [3]), .B(data[3]), .S(n_32), .Z(n_0_323));
   MUX2_X1 i_0_0_493 (.A(\mem[31] [2]), .B(data[2]), .S(n_32), .Z(n_0_322));
   MUX2_X1 i_0_0_494 (.A(\mem[31] [1]), .B(data[1]), .S(n_32), .Z(n_0_321));
   MUX2_X1 i_0_0_495 (.A(\mem[31] [0]), .B(data[0]), .S(n_32), .Z(n_0_320));
   MUX2_X1 i_0_0_496 (.A(\mem[32] [15]), .B(data[15]), .S(n_33), .Z(n_0_319));
   MUX2_X1 i_0_0_497 (.A(\mem[32] [14]), .B(data[14]), .S(n_33), .Z(n_0_318));
   MUX2_X1 i_0_0_498 (.A(\mem[32] [13]), .B(data[13]), .S(n_33), .Z(n_0_317));
   MUX2_X1 i_0_0_499 (.A(\mem[32] [12]), .B(data[12]), .S(n_33), .Z(n_0_316));
   MUX2_X1 i_0_0_500 (.A(\mem[32] [11]), .B(data[11]), .S(n_33), .Z(n_0_315));
   MUX2_X1 i_0_0_501 (.A(\mem[32] [10]), .B(data[10]), .S(n_33), .Z(n_0_314));
   MUX2_X1 i_0_0_502 (.A(\mem[32] [9]), .B(data[9]), .S(n_33), .Z(n_0_313));
   MUX2_X1 i_0_0_503 (.A(\mem[32] [8]), .B(data[8]), .S(n_33), .Z(n_0_312));
   MUX2_X1 i_0_0_504 (.A(\mem[32] [7]), .B(data[7]), .S(n_33), .Z(n_0_311));
   MUX2_X1 i_0_0_505 (.A(\mem[32] [6]), .B(data[6]), .S(n_33), .Z(n_0_310));
   MUX2_X1 i_0_0_506 (.A(\mem[32] [5]), .B(data[5]), .S(n_33), .Z(n_0_309));
   MUX2_X1 i_0_0_507 (.A(\mem[32] [4]), .B(data[4]), .S(n_33), .Z(n_0_308));
   MUX2_X1 i_0_0_508 (.A(\mem[32] [3]), .B(data[3]), .S(n_33), .Z(n_0_307));
   MUX2_X1 i_0_0_509 (.A(\mem[32] [2]), .B(data[2]), .S(n_33), .Z(n_0_306));
   MUX2_X1 i_0_0_510 (.A(\mem[32] [1]), .B(data[1]), .S(n_33), .Z(n_0_305));
   MUX2_X1 i_0_0_511 (.A(\mem[32] [0]), .B(data[0]), .S(n_33), .Z(n_0_304));
   MUX2_X1 i_0_0_512 (.A(\mem[33] [15]), .B(data[15]), .S(n_34), .Z(n_0_303));
   MUX2_X1 i_0_0_513 (.A(\mem[33] [14]), .B(data[14]), .S(n_34), .Z(n_0_302));
   MUX2_X1 i_0_0_514 (.A(\mem[33] [13]), .B(data[13]), .S(n_34), .Z(n_0_301));
   MUX2_X1 i_0_0_515 (.A(\mem[33] [12]), .B(data[12]), .S(n_34), .Z(n_0_300));
   MUX2_X1 i_0_0_516 (.A(\mem[33] [11]), .B(data[11]), .S(n_34), .Z(n_0_299));
   MUX2_X1 i_0_0_517 (.A(\mem[33] [10]), .B(data[10]), .S(n_34), .Z(n_0_298));
   MUX2_X1 i_0_0_518 (.A(\mem[33] [9]), .B(data[9]), .S(n_34), .Z(n_0_297));
   MUX2_X1 i_0_0_519 (.A(\mem[33] [8]), .B(data[8]), .S(n_34), .Z(n_0_296));
   MUX2_X1 i_0_0_520 (.A(\mem[33] [7]), .B(data[7]), .S(n_34), .Z(n_0_295));
   MUX2_X1 i_0_0_521 (.A(\mem[33] [6]), .B(data[6]), .S(n_34), .Z(n_0_294));
   MUX2_X1 i_0_0_522 (.A(\mem[33] [5]), .B(data[5]), .S(n_34), .Z(n_0_293));
   MUX2_X1 i_0_0_523 (.A(\mem[33] [4]), .B(data[4]), .S(n_34), .Z(n_0_292));
   MUX2_X1 i_0_0_524 (.A(\mem[33] [3]), .B(data[3]), .S(n_34), .Z(n_0_291));
   MUX2_X1 i_0_0_525 (.A(\mem[33] [2]), .B(data[2]), .S(n_34), .Z(n_0_290));
   MUX2_X1 i_0_0_526 (.A(\mem[33] [1]), .B(data[1]), .S(n_34), .Z(n_0_289));
   MUX2_X1 i_0_0_527 (.A(\mem[33] [0]), .B(data[0]), .S(n_34), .Z(n_0_288));
   MUX2_X1 i_0_0_528 (.A(\mem[34] [15]), .B(data[15]), .S(n_35), .Z(n_0_287));
   MUX2_X1 i_0_0_529 (.A(\mem[34] [14]), .B(data[14]), .S(n_35), .Z(n_0_286));
   MUX2_X1 i_0_0_530 (.A(\mem[34] [13]), .B(data[13]), .S(n_35), .Z(n_0_285));
   MUX2_X1 i_0_0_531 (.A(\mem[34] [12]), .B(data[12]), .S(n_35), .Z(n_0_284));
   MUX2_X1 i_0_0_532 (.A(\mem[34] [11]), .B(data[11]), .S(n_35), .Z(n_0_283));
   MUX2_X1 i_0_0_533 (.A(\mem[34] [10]), .B(data[10]), .S(n_35), .Z(n_0_282));
   MUX2_X1 i_0_0_534 (.A(\mem[34] [9]), .B(data[9]), .S(n_35), .Z(n_0_281));
   MUX2_X1 i_0_0_535 (.A(\mem[34] [8]), .B(data[8]), .S(n_35), .Z(n_0_280));
   MUX2_X1 i_0_0_536 (.A(\mem[34] [7]), .B(data[7]), .S(n_35), .Z(n_0_279));
   MUX2_X1 i_0_0_537 (.A(\mem[34] [6]), .B(data[6]), .S(n_35), .Z(n_0_278));
   MUX2_X1 i_0_0_538 (.A(\mem[34] [5]), .B(data[5]), .S(n_35), .Z(n_0_277));
   MUX2_X1 i_0_0_539 (.A(\mem[34] [4]), .B(data[4]), .S(n_35), .Z(n_0_276));
   MUX2_X1 i_0_0_540 (.A(\mem[34] [3]), .B(data[3]), .S(n_35), .Z(n_0_275));
   MUX2_X1 i_0_0_541 (.A(\mem[34] [2]), .B(data[2]), .S(n_35), .Z(n_0_274));
   MUX2_X1 i_0_0_542 (.A(\mem[34] [1]), .B(data[1]), .S(n_35), .Z(n_0_273));
   MUX2_X1 i_0_0_543 (.A(\mem[34] [0]), .B(data[0]), .S(n_35), .Z(n_0_272));
   MUX2_X1 i_0_0_544 (.A(\mem[35] [15]), .B(data[15]), .S(n_36), .Z(n_0_271));
   MUX2_X1 i_0_0_545 (.A(\mem[35] [14]), .B(data[14]), .S(n_36), .Z(n_0_270));
   MUX2_X1 i_0_0_546 (.A(\mem[35] [13]), .B(data[13]), .S(n_36), .Z(n_0_269));
   MUX2_X1 i_0_0_547 (.A(\mem[35] [12]), .B(data[12]), .S(n_36), .Z(n_0_268));
   MUX2_X1 i_0_0_548 (.A(\mem[35] [11]), .B(data[11]), .S(n_36), .Z(n_0_267));
   MUX2_X1 i_0_0_549 (.A(\mem[35] [10]), .B(data[10]), .S(n_36), .Z(n_0_266));
   MUX2_X1 i_0_0_550 (.A(\mem[35] [9]), .B(data[9]), .S(n_36), .Z(n_0_265));
   MUX2_X1 i_0_0_551 (.A(\mem[35] [8]), .B(data[8]), .S(n_36), .Z(n_0_264));
   MUX2_X1 i_0_0_552 (.A(\mem[35] [7]), .B(data[7]), .S(n_36), .Z(n_0_263));
   MUX2_X1 i_0_0_553 (.A(\mem[35] [6]), .B(data[6]), .S(n_36), .Z(n_0_262));
   MUX2_X1 i_0_0_554 (.A(\mem[35] [5]), .B(data[5]), .S(n_36), .Z(n_0_261));
   MUX2_X1 i_0_0_555 (.A(\mem[35] [4]), .B(data[4]), .S(n_36), .Z(n_0_260));
   MUX2_X1 i_0_0_556 (.A(\mem[35] [3]), .B(data[3]), .S(n_36), .Z(n_0_259));
   MUX2_X1 i_0_0_557 (.A(\mem[35] [2]), .B(data[2]), .S(n_36), .Z(n_0_258));
   MUX2_X1 i_0_0_558 (.A(\mem[35] [1]), .B(data[1]), .S(n_36), .Z(n_0_257));
   MUX2_X1 i_0_0_559 (.A(\mem[35] [0]), .B(data[0]), .S(n_36), .Z(n_0_256));
   MUX2_X1 i_0_0_560 (.A(\mem[36] [15]), .B(data[15]), .S(n_37), .Z(n_0_255));
   MUX2_X1 i_0_0_561 (.A(\mem[36] [14]), .B(data[14]), .S(n_37), .Z(n_0_254));
   MUX2_X1 i_0_0_562 (.A(\mem[36] [13]), .B(data[13]), .S(n_37), .Z(n_0_253));
   MUX2_X1 i_0_0_563 (.A(\mem[36] [12]), .B(data[12]), .S(n_37), .Z(n_0_252));
   MUX2_X1 i_0_0_564 (.A(\mem[36] [11]), .B(data[11]), .S(n_37), .Z(n_0_251));
   MUX2_X1 i_0_0_565 (.A(\mem[36] [10]), .B(data[10]), .S(n_37), .Z(n_0_250));
   MUX2_X1 i_0_0_566 (.A(\mem[36] [9]), .B(data[9]), .S(n_37), .Z(n_0_249));
   MUX2_X1 i_0_0_567 (.A(\mem[36] [8]), .B(data[8]), .S(n_37), .Z(n_0_248));
   MUX2_X1 i_0_0_568 (.A(\mem[36] [7]), .B(data[7]), .S(n_37), .Z(n_0_247));
   MUX2_X1 i_0_0_569 (.A(\mem[36] [6]), .B(data[6]), .S(n_37), .Z(n_0_246));
   MUX2_X1 i_0_0_570 (.A(\mem[36] [5]), .B(data[5]), .S(n_37), .Z(n_0_245));
   MUX2_X1 i_0_0_571 (.A(\mem[36] [4]), .B(data[4]), .S(n_37), .Z(n_0_244));
   MUX2_X1 i_0_0_572 (.A(\mem[36] [3]), .B(data[3]), .S(n_37), .Z(n_0_243));
   MUX2_X1 i_0_0_573 (.A(\mem[36] [2]), .B(data[2]), .S(n_37), .Z(n_0_242));
   MUX2_X1 i_0_0_574 (.A(\mem[36] [1]), .B(data[1]), .S(n_37), .Z(n_0_241));
   MUX2_X1 i_0_0_575 (.A(\mem[36] [0]), .B(data[0]), .S(n_37), .Z(n_0_240));
   MUX2_X1 i_0_0_576 (.A(\mem[37] [15]), .B(data[15]), .S(n_38), .Z(n_0_239));
   MUX2_X1 i_0_0_577 (.A(\mem[37] [14]), .B(data[14]), .S(n_38), .Z(n_0_238));
   MUX2_X1 i_0_0_578 (.A(\mem[37] [13]), .B(data[13]), .S(n_38), .Z(n_0_237));
   MUX2_X1 i_0_0_579 (.A(\mem[37] [12]), .B(data[12]), .S(n_38), .Z(n_0_236));
   MUX2_X1 i_0_0_580 (.A(\mem[37] [11]), .B(data[11]), .S(n_38), .Z(n_0_235));
   MUX2_X1 i_0_0_581 (.A(\mem[37] [10]), .B(data[10]), .S(n_38), .Z(n_0_234));
   MUX2_X1 i_0_0_582 (.A(\mem[37] [9]), .B(data[9]), .S(n_38), .Z(n_0_233));
   MUX2_X1 i_0_0_583 (.A(\mem[37] [8]), .B(data[8]), .S(n_38), .Z(n_0_232));
   MUX2_X1 i_0_0_584 (.A(\mem[37] [7]), .B(data[7]), .S(n_38), .Z(n_0_231));
   MUX2_X1 i_0_0_585 (.A(\mem[37] [6]), .B(data[6]), .S(n_38), .Z(n_0_230));
   MUX2_X1 i_0_0_586 (.A(\mem[37] [5]), .B(data[5]), .S(n_38), .Z(n_0_229));
   MUX2_X1 i_0_0_587 (.A(\mem[37] [4]), .B(data[4]), .S(n_38), .Z(n_0_228));
   MUX2_X1 i_0_0_588 (.A(\mem[37] [3]), .B(data[3]), .S(n_38), .Z(n_0_227));
   MUX2_X1 i_0_0_589 (.A(\mem[37] [2]), .B(data[2]), .S(n_38), .Z(n_0_226));
   MUX2_X1 i_0_0_590 (.A(\mem[37] [1]), .B(data[1]), .S(n_38), .Z(n_0_225));
   MUX2_X1 i_0_0_591 (.A(\mem[37] [0]), .B(data[0]), .S(n_38), .Z(n_0_224));
   MUX2_X1 i_0_0_592 (.A(\mem[38] [15]), .B(data[15]), .S(n_39), .Z(n_0_223));
   MUX2_X1 i_0_0_593 (.A(\mem[38] [14]), .B(data[14]), .S(n_39), .Z(n_0_222));
   MUX2_X1 i_0_0_594 (.A(\mem[38] [13]), .B(data[13]), .S(n_39), .Z(n_0_221));
   MUX2_X1 i_0_0_595 (.A(\mem[38] [12]), .B(data[12]), .S(n_39), .Z(n_0_220));
   MUX2_X1 i_0_0_596 (.A(\mem[38] [11]), .B(data[11]), .S(n_39), .Z(n_0_219));
   MUX2_X1 i_0_0_597 (.A(\mem[38] [10]), .B(data[10]), .S(n_39), .Z(n_0_218));
   MUX2_X1 i_0_0_598 (.A(\mem[38] [9]), .B(data[9]), .S(n_39), .Z(n_0_217));
   MUX2_X1 i_0_0_599 (.A(\mem[38] [8]), .B(data[8]), .S(n_39), .Z(n_0_216));
   MUX2_X1 i_0_0_600 (.A(\mem[38] [7]), .B(data[7]), .S(n_39), .Z(n_0_215));
   MUX2_X1 i_0_0_601 (.A(\mem[38] [6]), .B(data[6]), .S(n_39), .Z(n_0_214));
   MUX2_X1 i_0_0_602 (.A(\mem[38] [5]), .B(data[5]), .S(n_39), .Z(n_0_213));
   MUX2_X1 i_0_0_603 (.A(\mem[38] [4]), .B(data[4]), .S(n_39), .Z(n_0_212));
   MUX2_X1 i_0_0_604 (.A(\mem[38] [3]), .B(data[3]), .S(n_39), .Z(n_0_211));
   MUX2_X1 i_0_0_605 (.A(\mem[38] [2]), .B(data[2]), .S(n_39), .Z(n_0_210));
   MUX2_X1 i_0_0_606 (.A(\mem[38] [1]), .B(data[1]), .S(n_39), .Z(n_0_209));
   MUX2_X1 i_0_0_607 (.A(\mem[38] [0]), .B(data[0]), .S(n_39), .Z(n_0_208));
   MUX2_X1 i_0_0_608 (.A(\mem[39] [15]), .B(data[15]), .S(n_40), .Z(n_0_207));
   MUX2_X1 i_0_0_609 (.A(\mem[39] [14]), .B(data[14]), .S(n_40), .Z(n_0_206));
   MUX2_X1 i_0_0_610 (.A(\mem[39] [13]), .B(data[13]), .S(n_40), .Z(n_0_205));
   MUX2_X1 i_0_0_611 (.A(\mem[39] [12]), .B(data[12]), .S(n_40), .Z(n_0_204));
   MUX2_X1 i_0_0_612 (.A(\mem[39] [11]), .B(data[11]), .S(n_40), .Z(n_0_203));
   MUX2_X1 i_0_0_613 (.A(\mem[39] [10]), .B(data[10]), .S(n_40), .Z(n_0_202));
   MUX2_X1 i_0_0_614 (.A(\mem[39] [9]), .B(data[9]), .S(n_40), .Z(n_0_201));
   MUX2_X1 i_0_0_615 (.A(\mem[39] [8]), .B(data[8]), .S(n_40), .Z(n_0_200));
   MUX2_X1 i_0_0_616 (.A(\mem[39] [7]), .B(data[7]), .S(n_40), .Z(n_0_199));
   MUX2_X1 i_0_0_617 (.A(\mem[39] [6]), .B(data[6]), .S(n_40), .Z(n_0_198));
   MUX2_X1 i_0_0_618 (.A(\mem[39] [5]), .B(data[5]), .S(n_40), .Z(n_0_197));
   MUX2_X1 i_0_0_619 (.A(\mem[39] [4]), .B(data[4]), .S(n_40), .Z(n_0_196));
   MUX2_X1 i_0_0_620 (.A(\mem[39] [3]), .B(data[3]), .S(n_40), .Z(n_0_195));
   MUX2_X1 i_0_0_621 (.A(\mem[39] [2]), .B(data[2]), .S(n_40), .Z(n_0_194));
   MUX2_X1 i_0_0_622 (.A(\mem[39] [1]), .B(data[1]), .S(n_40), .Z(n_0_193));
   MUX2_X1 i_0_0_623 (.A(\mem[39] [0]), .B(data[0]), .S(n_40), .Z(n_0_192));
   MUX2_X1 i_0_0_624 (.A(\mem[40] [15]), .B(data[15]), .S(n_41), .Z(n_0_191));
   MUX2_X1 i_0_0_625 (.A(\mem[40] [14]), .B(data[14]), .S(n_41), .Z(n_0_190));
   MUX2_X1 i_0_0_626 (.A(\mem[40] [13]), .B(data[13]), .S(n_41), .Z(n_0_189));
   MUX2_X1 i_0_0_627 (.A(\mem[40] [12]), .B(data[12]), .S(n_41), .Z(n_0_188));
   MUX2_X1 i_0_0_628 (.A(\mem[40] [11]), .B(data[11]), .S(n_41), .Z(n_0_187));
   MUX2_X1 i_0_0_629 (.A(\mem[40] [10]), .B(data[10]), .S(n_41), .Z(n_0_186));
   MUX2_X1 i_0_0_630 (.A(\mem[40] [9]), .B(data[9]), .S(n_41), .Z(n_0_185));
   MUX2_X1 i_0_0_631 (.A(\mem[40] [8]), .B(data[8]), .S(n_41), .Z(n_0_184));
   MUX2_X1 i_0_0_632 (.A(\mem[40] [7]), .B(data[7]), .S(n_41), .Z(n_0_183));
   MUX2_X1 i_0_0_633 (.A(\mem[40] [6]), .B(data[6]), .S(n_41), .Z(n_0_182));
   MUX2_X1 i_0_0_634 (.A(\mem[40] [5]), .B(data[5]), .S(n_41), .Z(n_0_181));
   MUX2_X1 i_0_0_635 (.A(\mem[40] [4]), .B(data[4]), .S(n_41), .Z(n_0_180));
   MUX2_X1 i_0_0_636 (.A(\mem[40] [3]), .B(data[3]), .S(n_41), .Z(n_0_179));
   MUX2_X1 i_0_0_637 (.A(\mem[40] [2]), .B(data[2]), .S(n_41), .Z(n_0_178));
   MUX2_X1 i_0_0_638 (.A(\mem[40] [1]), .B(data[1]), .S(n_41), .Z(n_0_177));
   MUX2_X1 i_0_0_639 (.A(\mem[40] [0]), .B(data[0]), .S(n_41), .Z(n_0_176));
   MUX2_X1 i_0_0_640 (.A(\mem[41] [15]), .B(data[15]), .S(n_42), .Z(n_0_175));
   MUX2_X1 i_0_0_641 (.A(\mem[41] [14]), .B(data[14]), .S(n_42), .Z(n_0_174));
   MUX2_X1 i_0_0_642 (.A(\mem[41] [13]), .B(data[13]), .S(n_42), .Z(n_0_173));
   MUX2_X1 i_0_0_643 (.A(\mem[41] [12]), .B(data[12]), .S(n_42), .Z(n_0_172));
   MUX2_X1 i_0_0_644 (.A(\mem[41] [11]), .B(data[11]), .S(n_42), .Z(n_0_171));
   MUX2_X1 i_0_0_645 (.A(\mem[41] [10]), .B(data[10]), .S(n_42), .Z(n_0_170));
   MUX2_X1 i_0_0_646 (.A(\mem[41] [9]), .B(data[9]), .S(n_42), .Z(n_0_169));
   MUX2_X1 i_0_0_647 (.A(\mem[41] [8]), .B(data[8]), .S(n_42), .Z(n_0_168));
   MUX2_X1 i_0_0_648 (.A(\mem[41] [7]), .B(data[7]), .S(n_42), .Z(n_0_167));
   MUX2_X1 i_0_0_649 (.A(\mem[41] [6]), .B(data[6]), .S(n_42), .Z(n_0_166));
   MUX2_X1 i_0_0_650 (.A(\mem[41] [5]), .B(data[5]), .S(n_42), .Z(n_0_165));
   MUX2_X1 i_0_0_651 (.A(\mem[41] [4]), .B(data[4]), .S(n_42), .Z(n_0_164));
   MUX2_X1 i_0_0_652 (.A(\mem[41] [3]), .B(data[3]), .S(n_42), .Z(n_0_163));
   MUX2_X1 i_0_0_653 (.A(\mem[41] [2]), .B(data[2]), .S(n_42), .Z(n_0_162));
   MUX2_X1 i_0_0_654 (.A(\mem[41] [1]), .B(data[1]), .S(n_42), .Z(n_0_161));
   MUX2_X1 i_0_0_655 (.A(\mem[41] [0]), .B(data[0]), .S(n_42), .Z(n_0_160));
   MUX2_X1 i_0_0_656 (.A(\mem[42] [15]), .B(data[15]), .S(n_43), .Z(n_0_159));
   MUX2_X1 i_0_0_657 (.A(\mem[42] [14]), .B(data[14]), .S(n_43), .Z(n_0_158));
   MUX2_X1 i_0_0_658 (.A(\mem[42] [13]), .B(data[13]), .S(n_43), .Z(n_0_157));
   MUX2_X1 i_0_0_659 (.A(\mem[42] [12]), .B(data[12]), .S(n_43), .Z(n_0_156));
   MUX2_X1 i_0_0_660 (.A(\mem[42] [11]), .B(data[11]), .S(n_43), .Z(n_0_155));
   MUX2_X1 i_0_0_661 (.A(\mem[42] [10]), .B(data[10]), .S(n_43), .Z(n_0_154));
   MUX2_X1 i_0_0_662 (.A(\mem[42] [9]), .B(data[9]), .S(n_43), .Z(n_0_153));
   MUX2_X1 i_0_0_663 (.A(\mem[42] [8]), .B(data[8]), .S(n_43), .Z(n_0_152));
   MUX2_X1 i_0_0_664 (.A(\mem[42] [7]), .B(data[7]), .S(n_43), .Z(n_0_151));
   MUX2_X1 i_0_0_665 (.A(\mem[42] [6]), .B(data[6]), .S(n_43), .Z(n_0_150));
   MUX2_X1 i_0_0_666 (.A(\mem[42] [5]), .B(data[5]), .S(n_43), .Z(n_0_149));
   MUX2_X1 i_0_0_667 (.A(\mem[42] [4]), .B(data[4]), .S(n_43), .Z(n_0_148));
   MUX2_X1 i_0_0_668 (.A(\mem[42] [3]), .B(data[3]), .S(n_43), .Z(n_0_147));
   MUX2_X1 i_0_0_669 (.A(\mem[42] [2]), .B(data[2]), .S(n_43), .Z(n_0_146));
   MUX2_X1 i_0_0_670 (.A(\mem[42] [1]), .B(data[1]), .S(n_43), .Z(n_0_145));
   MUX2_X1 i_0_0_671 (.A(\mem[42] [0]), .B(data[0]), .S(n_43), .Z(n_0_144));
   MUX2_X1 i_0_0_672 (.A(\mem[43] [15]), .B(data[15]), .S(n_44), .Z(n_0_143));
   MUX2_X1 i_0_0_673 (.A(\mem[43] [14]), .B(data[14]), .S(n_44), .Z(n_0_142));
   MUX2_X1 i_0_0_674 (.A(\mem[43] [13]), .B(data[13]), .S(n_44), .Z(n_0_141));
   MUX2_X1 i_0_0_675 (.A(\mem[43] [12]), .B(data[12]), .S(n_44), .Z(n_0_140));
   MUX2_X1 i_0_0_676 (.A(\mem[43] [11]), .B(data[11]), .S(n_44), .Z(n_0_139));
   MUX2_X1 i_0_0_677 (.A(\mem[43] [10]), .B(data[10]), .S(n_44), .Z(n_0_138));
   MUX2_X1 i_0_0_678 (.A(\mem[43] [9]), .B(data[9]), .S(n_44), .Z(n_0_137));
   MUX2_X1 i_0_0_679 (.A(\mem[43] [8]), .B(data[8]), .S(n_44), .Z(n_0_136));
   MUX2_X1 i_0_0_680 (.A(\mem[43] [7]), .B(data[7]), .S(n_44), .Z(n_0_135));
   MUX2_X1 i_0_0_681 (.A(\mem[43] [6]), .B(data[6]), .S(n_44), .Z(n_0_134));
   MUX2_X1 i_0_0_682 (.A(\mem[43] [5]), .B(data[5]), .S(n_44), .Z(n_0_133));
   MUX2_X1 i_0_0_683 (.A(\mem[43] [4]), .B(data[4]), .S(n_44), .Z(n_0_132));
   MUX2_X1 i_0_0_684 (.A(\mem[43] [3]), .B(data[3]), .S(n_44), .Z(n_0_131));
   MUX2_X1 i_0_0_685 (.A(\mem[43] [2]), .B(data[2]), .S(n_44), .Z(n_0_130));
   MUX2_X1 i_0_0_686 (.A(\mem[43] [1]), .B(data[1]), .S(n_44), .Z(n_0_129));
   MUX2_X1 i_0_0_687 (.A(\mem[43] [0]), .B(data[0]), .S(n_44), .Z(n_0_128));
   MUX2_X1 i_0_0_688 (.A(\mem[44] [15]), .B(data[15]), .S(n_45), .Z(n_0_127));
   MUX2_X1 i_0_0_689 (.A(\mem[44] [14]), .B(data[14]), .S(n_45), .Z(n_0_126));
   MUX2_X1 i_0_0_690 (.A(\mem[44] [13]), .B(data[13]), .S(n_45), .Z(n_0_125));
   MUX2_X1 i_0_0_691 (.A(\mem[44] [12]), .B(data[12]), .S(n_45), .Z(n_0_124));
   MUX2_X1 i_0_0_692 (.A(\mem[44] [11]), .B(data[11]), .S(n_45), .Z(n_0_123));
   MUX2_X1 i_0_0_693 (.A(\mem[44] [10]), .B(data[10]), .S(n_45), .Z(n_0_122));
   MUX2_X1 i_0_0_694 (.A(\mem[44] [9]), .B(data[9]), .S(n_45), .Z(n_0_121));
   MUX2_X1 i_0_0_695 (.A(\mem[44] [8]), .B(data[8]), .S(n_45), .Z(n_0_120));
   MUX2_X1 i_0_0_696 (.A(\mem[44] [7]), .B(data[7]), .S(n_45), .Z(n_0_119));
   MUX2_X1 i_0_0_697 (.A(\mem[44] [6]), .B(data[6]), .S(n_45), .Z(n_0_118));
   MUX2_X1 i_0_0_698 (.A(\mem[44] [5]), .B(data[5]), .S(n_45), .Z(n_0_117));
   MUX2_X1 i_0_0_699 (.A(\mem[44] [4]), .B(data[4]), .S(n_45), .Z(n_0_116));
   MUX2_X1 i_0_0_700 (.A(\mem[44] [3]), .B(data[3]), .S(n_45), .Z(n_0_115));
   MUX2_X1 i_0_0_701 (.A(\mem[44] [2]), .B(data[2]), .S(n_45), .Z(n_0_114));
   MUX2_X1 i_0_0_702 (.A(\mem[44] [1]), .B(data[1]), .S(n_45), .Z(n_0_113));
   MUX2_X1 i_0_0_703 (.A(\mem[44] [0]), .B(data[0]), .S(n_45), .Z(n_0_112));
   MUX2_X1 i_0_0_704 (.A(\mem[45] [15]), .B(data[15]), .S(n_46), .Z(n_0_111));
   MUX2_X1 i_0_0_705 (.A(\mem[45] [14]), .B(data[14]), .S(n_46), .Z(n_0_110));
   MUX2_X1 i_0_0_706 (.A(\mem[45] [13]), .B(data[13]), .S(n_46), .Z(n_0_109));
   MUX2_X1 i_0_0_707 (.A(\mem[45] [12]), .B(data[12]), .S(n_46), .Z(n_0_108));
   MUX2_X1 i_0_0_708 (.A(\mem[45] [11]), .B(data[11]), .S(n_46), .Z(n_0_107));
   MUX2_X1 i_0_0_709 (.A(\mem[45] [10]), .B(data[10]), .S(n_46), .Z(n_0_106));
   MUX2_X1 i_0_0_710 (.A(\mem[45] [9]), .B(data[9]), .S(n_46), .Z(n_0_105));
   MUX2_X1 i_0_0_711 (.A(\mem[45] [8]), .B(data[8]), .S(n_46), .Z(n_0_104));
   MUX2_X1 i_0_0_712 (.A(\mem[45] [7]), .B(data[7]), .S(n_46), .Z(n_0_103));
   MUX2_X1 i_0_0_713 (.A(\mem[45] [6]), .B(data[6]), .S(n_46), .Z(n_0_102));
   MUX2_X1 i_0_0_714 (.A(\mem[45] [5]), .B(data[5]), .S(n_46), .Z(n_0_101));
   MUX2_X1 i_0_0_715 (.A(\mem[45] [4]), .B(data[4]), .S(n_46), .Z(n_0_100));
   MUX2_X1 i_0_0_716 (.A(\mem[45] [3]), .B(data[3]), .S(n_46), .Z(n_0_99));
   MUX2_X1 i_0_0_717 (.A(\mem[45] [2]), .B(data[2]), .S(n_46), .Z(n_0_98));
   MUX2_X1 i_0_0_718 (.A(\mem[45] [1]), .B(data[1]), .S(n_46), .Z(n_0_97));
   MUX2_X1 i_0_0_719 (.A(\mem[45] [0]), .B(data[0]), .S(n_46), .Z(n_0_96));
   MUX2_X1 i_0_0_720 (.A(\mem[46] [15]), .B(data[15]), .S(n_47), .Z(n_0_95));
   MUX2_X1 i_0_0_721 (.A(\mem[46] [14]), .B(data[14]), .S(n_47), .Z(n_0_94));
   MUX2_X1 i_0_0_722 (.A(\mem[46] [13]), .B(data[13]), .S(n_47), .Z(n_0_93));
   MUX2_X1 i_0_0_723 (.A(\mem[46] [12]), .B(data[12]), .S(n_47), .Z(n_0_92));
   MUX2_X1 i_0_0_724 (.A(\mem[46] [11]), .B(data[11]), .S(n_47), .Z(n_0_91));
   MUX2_X1 i_0_0_725 (.A(\mem[46] [10]), .B(data[10]), .S(n_47), .Z(n_0_90));
   MUX2_X1 i_0_0_726 (.A(\mem[46] [9]), .B(data[9]), .S(n_47), .Z(n_0_89));
   MUX2_X1 i_0_0_727 (.A(\mem[46] [8]), .B(data[8]), .S(n_47), .Z(n_0_88));
   MUX2_X1 i_0_0_728 (.A(\mem[46] [7]), .B(data[7]), .S(n_47), .Z(n_0_87));
   MUX2_X1 i_0_0_729 (.A(\mem[46] [6]), .B(data[6]), .S(n_47), .Z(n_0_86));
   MUX2_X1 i_0_0_730 (.A(\mem[46] [5]), .B(data[5]), .S(n_47), .Z(n_0_85));
   MUX2_X1 i_0_0_731 (.A(\mem[46] [4]), .B(data[4]), .S(n_47), .Z(n_0_84));
   MUX2_X1 i_0_0_732 (.A(\mem[46] [3]), .B(data[3]), .S(n_47), .Z(n_0_83));
   MUX2_X1 i_0_0_733 (.A(\mem[46] [2]), .B(data[2]), .S(n_47), .Z(n_0_82));
   MUX2_X1 i_0_0_734 (.A(\mem[46] [1]), .B(data[1]), .S(n_47), .Z(n_0_81));
   MUX2_X1 i_0_0_735 (.A(\mem[46] [0]), .B(data[0]), .S(n_47), .Z(n_0_80));
   MUX2_X1 i_0_0_736 (.A(\mem[47] [15]), .B(data[15]), .S(n_48), .Z(n_0_79));
   MUX2_X1 i_0_0_737 (.A(\mem[47] [14]), .B(data[14]), .S(n_48), .Z(n_0_78));
   MUX2_X1 i_0_0_738 (.A(\mem[47] [13]), .B(data[13]), .S(n_48), .Z(n_0_77));
   MUX2_X1 i_0_0_739 (.A(\mem[47] [12]), .B(data[12]), .S(n_48), .Z(n_0_76));
   MUX2_X1 i_0_0_740 (.A(\mem[47] [11]), .B(data[11]), .S(n_48), .Z(n_0_75));
   MUX2_X1 i_0_0_741 (.A(\mem[47] [10]), .B(data[10]), .S(n_48), .Z(n_0_74));
   MUX2_X1 i_0_0_742 (.A(\mem[47] [9]), .B(data[9]), .S(n_48), .Z(n_0_73));
   MUX2_X1 i_0_0_743 (.A(\mem[47] [8]), .B(data[8]), .S(n_48), .Z(n_0_72));
   MUX2_X1 i_0_0_744 (.A(\mem[47] [7]), .B(data[7]), .S(n_48), .Z(n_0_71));
   MUX2_X1 i_0_0_745 (.A(\mem[47] [6]), .B(data[6]), .S(n_48), .Z(n_0_70));
   MUX2_X1 i_0_0_746 (.A(\mem[47] [5]), .B(data[5]), .S(n_48), .Z(n_0_69));
   MUX2_X1 i_0_0_747 (.A(\mem[47] [4]), .B(data[4]), .S(n_48), .Z(n_0_68));
   MUX2_X1 i_0_0_748 (.A(\mem[47] [3]), .B(data[3]), .S(n_48), .Z(n_0_67));
   MUX2_X1 i_0_0_749 (.A(\mem[47] [2]), .B(data[2]), .S(n_48), .Z(n_0_66));
   MUX2_X1 i_0_0_750 (.A(\mem[47] [1]), .B(data[1]), .S(n_48), .Z(n_0_65));
   MUX2_X1 i_0_0_751 (.A(\mem[47] [0]), .B(data[0]), .S(n_48), .Z(n_0_64));
   MUX2_X1 i_0_0_752 (.A(\mem[48] [15]), .B(data[15]), .S(n_49), .Z(n_0_63));
   MUX2_X1 i_0_0_753 (.A(\mem[48] [14]), .B(data[14]), .S(n_49), .Z(n_0_62));
   MUX2_X1 i_0_0_754 (.A(\mem[48] [13]), .B(data[13]), .S(n_49), .Z(n_0_61));
   MUX2_X1 i_0_0_755 (.A(\mem[48] [12]), .B(data[12]), .S(n_49), .Z(n_0_60));
   MUX2_X1 i_0_0_756 (.A(\mem[48] [11]), .B(data[11]), .S(n_49), .Z(n_0_59));
   MUX2_X1 i_0_0_757 (.A(\mem[48] [10]), .B(data[10]), .S(n_49), .Z(n_0_58));
   MUX2_X1 i_0_0_758 (.A(\mem[48] [9]), .B(data[9]), .S(n_49), .Z(n_0_57));
   MUX2_X1 i_0_0_759 (.A(\mem[48] [8]), .B(data[8]), .S(n_49), .Z(n_0_56));
   MUX2_X1 i_0_0_760 (.A(\mem[48] [7]), .B(data[7]), .S(n_49), .Z(n_0_55));
   MUX2_X1 i_0_0_761 (.A(\mem[48] [6]), .B(data[6]), .S(n_49), .Z(n_0_54));
   MUX2_X1 i_0_0_762 (.A(\mem[48] [5]), .B(data[5]), .S(n_49), .Z(n_0_53));
   MUX2_X1 i_0_0_763 (.A(\mem[48] [4]), .B(data[4]), .S(n_49), .Z(n_0_52));
   MUX2_X1 i_0_0_764 (.A(\mem[48] [3]), .B(data[3]), .S(n_49), .Z(n_0_51));
   MUX2_X1 i_0_0_765 (.A(\mem[48] [2]), .B(data[2]), .S(n_49), .Z(n_0_50));
   MUX2_X1 i_0_0_766 (.A(\mem[48] [1]), .B(data[1]), .S(n_49), .Z(n_0_49));
   MUX2_X1 i_0_0_767 (.A(\mem[48] [0]), .B(data[0]), .S(n_49), .Z(n_0_48));
   MUX2_X1 i_0_0_768 (.A(\mem[49] [15]), .B(data[15]), .S(n_50), .Z(n_0_47));
   MUX2_X1 i_0_0_769 (.A(\mem[49] [14]), .B(data[14]), .S(n_50), .Z(n_0_46));
   MUX2_X1 i_0_0_770 (.A(\mem[49] [13]), .B(data[13]), .S(n_50), .Z(n_0_45));
   MUX2_X1 i_0_0_771 (.A(\mem[49] [12]), .B(data[12]), .S(n_50), .Z(n_0_44));
   MUX2_X1 i_0_0_772 (.A(\mem[49] [11]), .B(data[11]), .S(n_50), .Z(n_0_43));
   MUX2_X1 i_0_0_773 (.A(\mem[49] [10]), .B(data[10]), .S(n_50), .Z(n_0_42));
   MUX2_X1 i_0_0_774 (.A(\mem[49] [9]), .B(data[9]), .S(n_50), .Z(n_0_41));
   MUX2_X1 i_0_0_775 (.A(\mem[49] [8]), .B(data[8]), .S(n_50), .Z(n_0_40));
   MUX2_X1 i_0_0_776 (.A(\mem[49] [7]), .B(data[7]), .S(n_50), .Z(n_0_39));
   MUX2_X1 i_0_0_777 (.A(\mem[49] [6]), .B(data[6]), .S(n_50), .Z(n_0_38));
   MUX2_X1 i_0_0_778 (.A(\mem[49] [5]), .B(data[5]), .S(n_50), .Z(n_0_37));
   MUX2_X1 i_0_0_779 (.A(\mem[49] [4]), .B(data[4]), .S(n_50), .Z(n_0_36));
   MUX2_X1 i_0_0_780 (.A(\mem[49] [3]), .B(data[3]), .S(n_50), .Z(n_0_35));
   MUX2_X1 i_0_0_781 (.A(\mem[49] [2]), .B(data[2]), .S(n_50), .Z(n_0_34));
   MUX2_X1 i_0_0_782 (.A(\mem[49] [1]), .B(data[1]), .S(n_50), .Z(n_0_33));
   MUX2_X1 i_0_0_783 (.A(\mem[49] [0]), .B(data[0]), .S(n_50), .Z(n_0_32));
   MUX2_X1 i_0_0_784 (.A(\mem[51] [15]), .B(data[15]), .S(n_52), .Z(n_0_31));
   MUX2_X1 i_0_0_785 (.A(\mem[51] [14]), .B(data[14]), .S(n_52), .Z(n_0_30));
   MUX2_X1 i_0_0_786 (.A(\mem[51] [13]), .B(data[13]), .S(n_52), .Z(n_0_29));
   MUX2_X1 i_0_0_787 (.A(\mem[51] [12]), .B(data[12]), .S(n_52), .Z(n_0_28));
   MUX2_X1 i_0_0_788 (.A(\mem[51] [11]), .B(data[11]), .S(n_52), .Z(n_0_27));
   MUX2_X1 i_0_0_789 (.A(\mem[51] [10]), .B(data[10]), .S(n_52), .Z(n_0_26));
   MUX2_X1 i_0_0_790 (.A(\mem[51] [9]), .B(data[9]), .S(n_52), .Z(n_0_25));
   MUX2_X1 i_0_0_791 (.A(\mem[51] [8]), .B(data[8]), .S(n_52), .Z(n_0_24));
   MUX2_X1 i_0_0_792 (.A(\mem[51] [7]), .B(data[7]), .S(n_52), .Z(n_0_23));
   MUX2_X1 i_0_0_793 (.A(\mem[51] [6]), .B(data[6]), .S(n_52), .Z(n_0_22));
   MUX2_X1 i_0_0_794 (.A(\mem[51] [5]), .B(data[5]), .S(n_52), .Z(n_0_21));
   MUX2_X1 i_0_0_795 (.A(\mem[51] [4]), .B(data[4]), .S(n_52), .Z(n_0_20));
   MUX2_X1 i_0_0_796 (.A(\mem[51] [3]), .B(data[3]), .S(n_52), .Z(n_0_19));
   MUX2_X1 i_0_0_797 (.A(\mem[51] [2]), .B(data[2]), .S(n_52), .Z(n_0_18));
   MUX2_X1 i_0_0_798 (.A(\mem[51] [1]), .B(data[1]), .S(n_52), .Z(n_0_17));
   MUX2_X1 i_0_0_799 (.A(\mem[51] [0]), .B(data[0]), .S(n_52), .Z(n_0_16));
   MUX2_X1 i_0_0_800 (.A(\mem[50] [15]), .B(data[15]), .S(n_51), .Z(n_0_15));
   MUX2_X1 i_0_0_801 (.A(\mem[50] [14]), .B(data[14]), .S(n_51), .Z(n_0_14));
   MUX2_X1 i_0_0_802 (.A(\mem[50] [13]), .B(data[13]), .S(n_51), .Z(n_0_13));
   MUX2_X1 i_0_0_803 (.A(\mem[50] [12]), .B(data[12]), .S(n_51), .Z(n_0_12));
   MUX2_X1 i_0_0_804 (.A(\mem[50] [11]), .B(data[11]), .S(n_51), .Z(n_0_11));
   MUX2_X1 i_0_0_805 (.A(\mem[50] [10]), .B(data[10]), .S(n_51), .Z(n_0_10));
   MUX2_X1 i_0_0_806 (.A(\mem[50] [9]), .B(data[9]), .S(n_51), .Z(n_0_9));
   MUX2_X1 i_0_0_807 (.A(\mem[50] [8]), .B(data[8]), .S(n_51), .Z(n_0_8));
   MUX2_X1 i_0_0_808 (.A(\mem[50] [7]), .B(data[7]), .S(n_51), .Z(n_0_7));
   MUX2_X1 i_0_0_809 (.A(\mem[50] [6]), .B(data[6]), .S(n_51), .Z(n_0_6));
   MUX2_X1 i_0_0_810 (.A(\mem[50] [5]), .B(data[5]), .S(n_51), .Z(n_0_5));
   MUX2_X1 i_0_0_811 (.A(\mem[50] [4]), .B(data[4]), .S(n_51), .Z(n_0_4));
   MUX2_X1 i_0_0_812 (.A(\mem[50] [3]), .B(data[3]), .S(n_51), .Z(n_0_3));
   MUX2_X1 i_0_0_813 (.A(\mem[50] [2]), .B(data[2]), .S(n_51), .Z(n_0_2));
   MUX2_X1 i_0_0_814 (.A(\mem[50] [1]), .B(data[1]), .S(n_51), .Z(n_0_1));
   MUX2_X1 i_0_0_815 (.A(\mem[50] [0]), .B(data[0]), .S(n_51), .Z(n_0_0));
   DFF_X1 \mem_reg[52][15]  (.D(n_106_799), .CK(n_0), .Q(\mem[52] [15]), .QN());
   DFF_X1 \mem_reg[52][14]  (.D(n_106_798), .CK(n_0), .Q(\mem[52] [14]), .QN());
   DFF_X1 \mem_reg[52][13]  (.D(n_106_797), .CK(n_0), .Q(\mem[52] [13]), .QN());
   DFF_X1 \mem_reg[52][12]  (.D(n_106_796), .CK(n_0), .Q(\mem[52] [12]), .QN());
   DFF_X1 \mem_reg[52][11]  (.D(n_106_795), .CK(n_0), .Q(\mem[52] [11]), .QN());
   DFF_X1 \mem_reg[52][10]  (.D(n_106_794), .CK(n_0), .Q(\mem[52] [10]), .QN());
   DFF_X1 \mem_reg[52][9]  (.D(n_106_793), .CK(n_0), .Q(\mem[52] [9]), .QN());
   DFF_X1 \mem_reg[52][8]  (.D(n_106_792), .CK(n_0), .Q(\mem[52] [8]), .QN());
   DFF_X1 \mem_reg[52][7]  (.D(n_106_791), .CK(n_0), .Q(\mem[52] [7]), .QN());
   DFF_X1 \mem_reg[52][6]  (.D(n_106_790), .CK(n_0), .Q(\mem[52] [6]), .QN());
   DFF_X1 \mem_reg[52][5]  (.D(n_106_789), .CK(n_0), .Q(\mem[52] [5]), .QN());
   DFF_X1 \mem_reg[52][4]  (.D(n_106_788), .CK(n_0), .Q(\mem[52] [4]), .QN());
   DFF_X1 \mem_reg[52][3]  (.D(n_106_787), .CK(n_0), .Q(\mem[52] [3]), .QN());
   DFF_X1 \mem_reg[52][2]  (.D(n_106_786), .CK(n_0), .Q(\mem[52] [2]), .QN());
   DFF_X1 \mem_reg[52][1]  (.D(n_106_785), .CK(n_0), .Q(\mem[52] [1]), .QN());
   DFF_X1 \mem_reg[52][0]  (.D(n_106_784), .CK(n_0), .Q(\mem[52] [0]), .QN());
   DFF_X1 \mem_reg[53][15]  (.D(n_106_783), .CK(n_0), .Q(\mem[53] [15]), .QN());
   DFF_X1 \mem_reg[53][14]  (.D(n_106_782), .CK(n_0), .Q(\mem[53] [14]), .QN());
   DFF_X1 \mem_reg[53][13]  (.D(n_106_781), .CK(n_0), .Q(\mem[53] [13]), .QN());
   DFF_X1 \mem_reg[53][12]  (.D(n_106_780), .CK(n_0), .Q(\mem[53] [12]), .QN());
   DFF_X1 \mem_reg[53][11]  (.D(n_106_779), .CK(n_0), .Q(\mem[53] [11]), .QN());
   DFF_X1 \mem_reg[53][10]  (.D(n_106_778), .CK(n_0), .Q(\mem[53] [10]), .QN());
   DFF_X1 \mem_reg[53][9]  (.D(n_106_777), .CK(n_0), .Q(\mem[53] [9]), .QN());
   DFF_X1 \mem_reg[53][8]  (.D(n_106_776), .CK(n_0), .Q(\mem[53] [8]), .QN());
   DFF_X1 \mem_reg[53][7]  (.D(n_106_775), .CK(n_0), .Q(\mem[53] [7]), .QN());
   DFF_X1 \mem_reg[53][6]  (.D(n_106_774), .CK(n_0), .Q(\mem[53] [6]), .QN());
   DFF_X1 \mem_reg[53][5]  (.D(n_106_773), .CK(n_0), .Q(\mem[53] [5]), .QN());
   DFF_X1 \mem_reg[53][4]  (.D(n_106_772), .CK(n_0), .Q(\mem[53] [4]), .QN());
   DFF_X1 \mem_reg[53][3]  (.D(n_106_771), .CK(n_0), .Q(\mem[53] [3]), .QN());
   DFF_X1 \mem_reg[53][2]  (.D(n_106_770), .CK(n_0), .Q(\mem[53] [2]), .QN());
   DFF_X1 \mem_reg[53][1]  (.D(n_106_769), .CK(n_0), .Q(\mem[53] [1]), .QN());
   DFF_X1 \mem_reg[53][0]  (.D(n_106_768), .CK(n_0), .Q(\mem[53] [0]), .QN());
   DFF_X1 \mem_reg[54][15]  (.D(n_106_767), .CK(n_0), .Q(\mem[54] [15]), .QN());
   DFF_X1 \mem_reg[54][14]  (.D(n_106_766), .CK(n_0), .Q(\mem[54] [14]), .QN());
   DFF_X1 \mem_reg[54][13]  (.D(n_106_765), .CK(n_0), .Q(\mem[54] [13]), .QN());
   DFF_X1 \mem_reg[54][12]  (.D(n_106_764), .CK(n_0), .Q(\mem[54] [12]), .QN());
   DFF_X1 \mem_reg[54][11]  (.D(n_106_763), .CK(n_0), .Q(\mem[54] [11]), .QN());
   DFF_X1 \mem_reg[54][10]  (.D(n_106_762), .CK(n_0), .Q(\mem[54] [10]), .QN());
   DFF_X1 \mem_reg[54][9]  (.D(n_106_761), .CK(n_0), .Q(\mem[54] [9]), .QN());
   DFF_X1 \mem_reg[54][8]  (.D(n_106_760), .CK(n_0), .Q(\mem[54] [8]), .QN());
   DFF_X1 \mem_reg[54][7]  (.D(n_106_759), .CK(n_0), .Q(\mem[54] [7]), .QN());
   DFF_X1 \mem_reg[54][6]  (.D(n_106_758), .CK(n_0), .Q(\mem[54] [6]), .QN());
   DFF_X1 \mem_reg[54][5]  (.D(n_106_757), .CK(n_0), .Q(\mem[54] [5]), .QN());
   DFF_X1 \mem_reg[54][4]  (.D(n_106_756), .CK(n_0), .Q(\mem[54] [4]), .QN());
   DFF_X1 \mem_reg[54][3]  (.D(n_106_755), .CK(n_0), .Q(\mem[54] [3]), .QN());
   DFF_X1 \mem_reg[54][2]  (.D(n_106_754), .CK(n_0), .Q(\mem[54] [2]), .QN());
   DFF_X1 \mem_reg[54][1]  (.D(n_106_753), .CK(n_0), .Q(\mem[54] [1]), .QN());
   DFF_X1 \mem_reg[54][0]  (.D(n_106_752), .CK(n_0), .Q(\mem[54] [0]), .QN());
   DFF_X1 \mem_reg[55][15]  (.D(n_106_751), .CK(n_0), .Q(\mem[55] [15]), .QN());
   DFF_X1 \mem_reg[55][14]  (.D(n_106_750), .CK(n_0), .Q(\mem[55] [14]), .QN());
   DFF_X1 \mem_reg[55][13]  (.D(n_106_749), .CK(n_0), .Q(\mem[55] [13]), .QN());
   DFF_X1 \mem_reg[55][12]  (.D(n_106_748), .CK(n_0), .Q(\mem[55] [12]), .QN());
   DFF_X1 \mem_reg[55][11]  (.D(n_106_747), .CK(n_0), .Q(\mem[55] [11]), .QN());
   DFF_X1 \mem_reg[55][10]  (.D(n_106_746), .CK(n_0), .Q(\mem[55] [10]), .QN());
   DFF_X1 \mem_reg[55][9]  (.D(n_106_745), .CK(n_0), .Q(\mem[55] [9]), .QN());
   DFF_X1 \mem_reg[55][8]  (.D(n_106_744), .CK(n_0), .Q(\mem[55] [8]), .QN());
   DFF_X1 \mem_reg[55][7]  (.D(n_106_743), .CK(n_0), .Q(\mem[55] [7]), .QN());
   DFF_X1 \mem_reg[55][6]  (.D(n_106_742), .CK(n_0), .Q(\mem[55] [6]), .QN());
   DFF_X1 \mem_reg[55][5]  (.D(n_106_741), .CK(n_0), .Q(\mem[55] [5]), .QN());
   DFF_X1 \mem_reg[55][4]  (.D(n_106_740), .CK(n_0), .Q(\mem[55] [4]), .QN());
   DFF_X1 \mem_reg[55][3]  (.D(n_106_739), .CK(n_0), .Q(\mem[55] [3]), .QN());
   DFF_X1 \mem_reg[55][2]  (.D(n_106_738), .CK(n_0), .Q(\mem[55] [2]), .QN());
   DFF_X1 \mem_reg[55][1]  (.D(n_106_737), .CK(n_0), .Q(\mem[55] [1]), .QN());
   DFF_X1 \mem_reg[55][0]  (.D(n_106_736), .CK(n_0), .Q(\mem[55] [0]), .QN());
   DFF_X1 \mem_reg[56][15]  (.D(n_106_735), .CK(n_0), .Q(\mem[56] [15]), .QN());
   DFF_X1 \mem_reg[56][14]  (.D(n_106_734), .CK(n_0), .Q(\mem[56] [14]), .QN());
   DFF_X1 \mem_reg[56][13]  (.D(n_106_733), .CK(n_0), .Q(\mem[56] [13]), .QN());
   DFF_X1 \mem_reg[56][12]  (.D(n_106_732), .CK(n_0), .Q(\mem[56] [12]), .QN());
   DFF_X1 \mem_reg[56][11]  (.D(n_106_731), .CK(n_0), .Q(\mem[56] [11]), .QN());
   DFF_X1 \mem_reg[56][10]  (.D(n_106_730), .CK(n_0), .Q(\mem[56] [10]), .QN());
   DFF_X1 \mem_reg[56][9]  (.D(n_106_729), .CK(n_0), .Q(\mem[56] [9]), .QN());
   DFF_X1 \mem_reg[56][8]  (.D(n_106_728), .CK(n_0), .Q(\mem[56] [8]), .QN());
   DFF_X1 \mem_reg[56][7]  (.D(n_106_727), .CK(n_0), .Q(\mem[56] [7]), .QN());
   DFF_X1 \mem_reg[56][6]  (.D(n_106_726), .CK(n_0), .Q(\mem[56] [6]), .QN());
   DFF_X1 \mem_reg[56][5]  (.D(n_106_725), .CK(n_0), .Q(\mem[56] [5]), .QN());
   DFF_X1 \mem_reg[56][4]  (.D(n_106_724), .CK(n_0), .Q(\mem[56] [4]), .QN());
   DFF_X1 \mem_reg[56][3]  (.D(n_106_723), .CK(n_0), .Q(\mem[56] [3]), .QN());
   DFF_X1 \mem_reg[56][2]  (.D(n_106_722), .CK(n_0), .Q(\mem[56] [2]), .QN());
   DFF_X1 \mem_reg[56][1]  (.D(n_106_721), .CK(n_0), .Q(\mem[56] [1]), .QN());
   DFF_X1 \mem_reg[56][0]  (.D(n_106_720), .CK(n_0), .Q(\mem[56] [0]), .QN());
   DFF_X1 \mem_reg[57][15]  (.D(n_106_719), .CK(n_0), .Q(\mem[57] [15]), .QN());
   DFF_X1 \mem_reg[57][14]  (.D(n_106_718), .CK(n_0), .Q(\mem[57] [14]), .QN());
   DFF_X1 \mem_reg[57][13]  (.D(n_106_717), .CK(n_0), .Q(\mem[57] [13]), .QN());
   DFF_X1 \mem_reg[57][12]  (.D(n_106_716), .CK(n_0), .Q(\mem[57] [12]), .QN());
   DFF_X1 \mem_reg[57][11]  (.D(n_106_715), .CK(n_0), .Q(\mem[57] [11]), .QN());
   DFF_X1 \mem_reg[57][10]  (.D(n_106_714), .CK(n_0), .Q(\mem[57] [10]), .QN());
   DFF_X1 \mem_reg[57][9]  (.D(n_106_713), .CK(n_0), .Q(\mem[57] [9]), .QN());
   DFF_X1 \mem_reg[57][8]  (.D(n_106_712), .CK(n_0), .Q(\mem[57] [8]), .QN());
   DFF_X1 \mem_reg[57][7]  (.D(n_106_711), .CK(n_0), .Q(\mem[57] [7]), .QN());
   DFF_X1 \mem_reg[57][6]  (.D(n_106_710), .CK(n_0), .Q(\mem[57] [6]), .QN());
   DFF_X1 \mem_reg[57][5]  (.D(n_106_709), .CK(n_0), .Q(\mem[57] [5]), .QN());
   DFF_X1 \mem_reg[57][4]  (.D(n_106_708), .CK(n_0), .Q(\mem[57] [4]), .QN());
   DFF_X1 \mem_reg[57][3]  (.D(n_106_707), .CK(n_0), .Q(\mem[57] [3]), .QN());
   DFF_X1 \mem_reg[57][2]  (.D(n_106_706), .CK(n_0), .Q(\mem[57] [2]), .QN());
   DFF_X1 \mem_reg[57][1]  (.D(n_106_705), .CK(n_0), .Q(\mem[57] [1]), .QN());
   DFF_X1 \mem_reg[57][0]  (.D(n_106_704), .CK(n_0), .Q(\mem[57] [0]), .QN());
   DFF_X1 \mem_reg[58][15]  (.D(n_106_703), .CK(n_0), .Q(\mem[58] [15]), .QN());
   DFF_X1 \mem_reg[58][14]  (.D(n_106_702), .CK(n_0), .Q(\mem[58] [14]), .QN());
   DFF_X1 \mem_reg[58][13]  (.D(n_106_701), .CK(n_0), .Q(\mem[58] [13]), .QN());
   DFF_X1 \mem_reg[58][12]  (.D(n_106_700), .CK(n_0), .Q(\mem[58] [12]), .QN());
   DFF_X1 \mem_reg[58][11]  (.D(n_106_699), .CK(n_0), .Q(\mem[58] [11]), .QN());
   DFF_X1 \mem_reg[58][10]  (.D(n_106_698), .CK(n_0), .Q(\mem[58] [10]), .QN());
   DFF_X1 \mem_reg[58][9]  (.D(n_106_697), .CK(n_0), .Q(\mem[58] [9]), .QN());
   DFF_X1 \mem_reg[58][8]  (.D(n_106_696), .CK(n_0), .Q(\mem[58] [8]), .QN());
   DFF_X1 \mem_reg[58][7]  (.D(n_106_695), .CK(n_0), .Q(\mem[58] [7]), .QN());
   DFF_X1 \mem_reg[58][6]  (.D(n_106_694), .CK(n_0), .Q(\mem[58] [6]), .QN());
   DFF_X1 \mem_reg[58][5]  (.D(n_106_693), .CK(n_0), .Q(\mem[58] [5]), .QN());
   DFF_X1 \mem_reg[58][4]  (.D(n_106_692), .CK(n_0), .Q(\mem[58] [4]), .QN());
   DFF_X1 \mem_reg[58][3]  (.D(n_106_691), .CK(n_0), .Q(\mem[58] [3]), .QN());
   DFF_X1 \mem_reg[58][2]  (.D(n_106_690), .CK(n_0), .Q(\mem[58] [2]), .QN());
   DFF_X1 \mem_reg[58][1]  (.D(n_106_689), .CK(n_0), .Q(\mem[58] [1]), .QN());
   DFF_X1 \mem_reg[58][0]  (.D(n_106_688), .CK(n_0), .Q(\mem[58] [0]), .QN());
   DFF_X1 \mem_reg[59][15]  (.D(n_106_687), .CK(n_0), .Q(\mem[59] [15]), .QN());
   DFF_X1 \mem_reg[59][14]  (.D(n_106_686), .CK(n_0), .Q(\mem[59] [14]), .QN());
   DFF_X1 \mem_reg[59][13]  (.D(n_106_685), .CK(n_0), .Q(\mem[59] [13]), .QN());
   DFF_X1 \mem_reg[59][12]  (.D(n_106_684), .CK(n_0), .Q(\mem[59] [12]), .QN());
   DFF_X1 \mem_reg[59][11]  (.D(n_106_683), .CK(n_0), .Q(\mem[59] [11]), .QN());
   DFF_X1 \mem_reg[59][10]  (.D(n_106_682), .CK(n_0), .Q(\mem[59] [10]), .QN());
   DFF_X1 \mem_reg[59][9]  (.D(n_106_681), .CK(n_0), .Q(\mem[59] [9]), .QN());
   DFF_X1 \mem_reg[59][8]  (.D(n_106_680), .CK(n_0), .Q(\mem[59] [8]), .QN());
   DFF_X1 \mem_reg[59][7]  (.D(n_106_679), .CK(n_0), .Q(\mem[59] [7]), .QN());
   DFF_X1 \mem_reg[59][6]  (.D(n_106_678), .CK(n_0), .Q(\mem[59] [6]), .QN());
   DFF_X1 \mem_reg[59][5]  (.D(n_106_677), .CK(n_0), .Q(\mem[59] [5]), .QN());
   DFF_X1 \mem_reg[59][4]  (.D(n_106_676), .CK(n_0), .Q(\mem[59] [4]), .QN());
   DFF_X1 \mem_reg[59][3]  (.D(n_106_675), .CK(n_0), .Q(\mem[59] [3]), .QN());
   DFF_X1 \mem_reg[59][2]  (.D(n_106_674), .CK(n_0), .Q(\mem[59] [2]), .QN());
   DFF_X1 \mem_reg[59][1]  (.D(n_106_673), .CK(n_0), .Q(\mem[59] [1]), .QN());
   DFF_X1 \mem_reg[59][0]  (.D(n_106_672), .CK(n_0), .Q(\mem[59] [0]), .QN());
   DFF_X1 \mem_reg[60][15]  (.D(n_106_671), .CK(n_0), .Q(\mem[60] [15]), .QN());
   DFF_X1 \mem_reg[60][14]  (.D(n_106_670), .CK(n_0), .Q(\mem[60] [14]), .QN());
   DFF_X1 \mem_reg[60][13]  (.D(n_106_669), .CK(n_0), .Q(\mem[60] [13]), .QN());
   DFF_X1 \mem_reg[60][12]  (.D(n_106_668), .CK(n_0), .Q(\mem[60] [12]), .QN());
   DFF_X1 \mem_reg[60][11]  (.D(n_106_667), .CK(n_0), .Q(\mem[60] [11]), .QN());
   DFF_X1 \mem_reg[60][10]  (.D(n_106_666), .CK(n_0), .Q(\mem[60] [10]), .QN());
   DFF_X1 \mem_reg[60][9]  (.D(n_106_665), .CK(n_0), .Q(\mem[60] [9]), .QN());
   DFF_X1 \mem_reg[60][8]  (.D(n_106_664), .CK(n_0), .Q(\mem[60] [8]), .QN());
   DFF_X1 \mem_reg[60][7]  (.D(n_106_663), .CK(n_0), .Q(\mem[60] [7]), .QN());
   DFF_X1 \mem_reg[60][6]  (.D(n_106_662), .CK(n_0), .Q(\mem[60] [6]), .QN());
   DFF_X1 \mem_reg[60][5]  (.D(n_106_661), .CK(n_0), .Q(\mem[60] [5]), .QN());
   DFF_X1 \mem_reg[60][4]  (.D(n_106_660), .CK(n_0), .Q(\mem[60] [4]), .QN());
   DFF_X1 \mem_reg[60][3]  (.D(n_106_659), .CK(n_0), .Q(\mem[60] [3]), .QN());
   DFF_X1 \mem_reg[60][2]  (.D(n_106_658), .CK(n_0), .Q(\mem[60] [2]), .QN());
   DFF_X1 \mem_reg[60][1]  (.D(n_106_657), .CK(n_0), .Q(\mem[60] [1]), .QN());
   DFF_X1 \mem_reg[60][0]  (.D(n_106_656), .CK(n_0), .Q(\mem[60] [0]), .QN());
   DFF_X1 \mem_reg[61][15]  (.D(n_106_655), .CK(n_0), .Q(\mem[61] [15]), .QN());
   DFF_X1 \mem_reg[61][14]  (.D(n_106_654), .CK(n_0), .Q(\mem[61] [14]), .QN());
   DFF_X1 \mem_reg[61][13]  (.D(n_106_653), .CK(n_0), .Q(\mem[61] [13]), .QN());
   DFF_X1 \mem_reg[61][12]  (.D(n_106_652), .CK(n_0), .Q(\mem[61] [12]), .QN());
   DFF_X1 \mem_reg[61][11]  (.D(n_106_651), .CK(n_0), .Q(\mem[61] [11]), .QN());
   DFF_X1 \mem_reg[61][10]  (.D(n_106_650), .CK(n_0), .Q(\mem[61] [10]), .QN());
   DFF_X1 \mem_reg[61][9]  (.D(n_106_649), .CK(n_0), .Q(\mem[61] [9]), .QN());
   DFF_X1 \mem_reg[61][8]  (.D(n_106_648), .CK(n_0), .Q(\mem[61] [8]), .QN());
   DFF_X1 \mem_reg[61][7]  (.D(n_106_647), .CK(n_0), .Q(\mem[61] [7]), .QN());
   DFF_X1 \mem_reg[61][6]  (.D(n_106_646), .CK(n_0), .Q(\mem[61] [6]), .QN());
   DFF_X1 \mem_reg[61][5]  (.D(n_106_645), .CK(n_0), .Q(\mem[61] [5]), .QN());
   DFF_X1 \mem_reg[61][4]  (.D(n_106_644), .CK(n_0), .Q(\mem[61] [4]), .QN());
   DFF_X1 \mem_reg[61][3]  (.D(n_106_643), .CK(n_0), .Q(\mem[61] [3]), .QN());
   DFF_X1 \mem_reg[61][2]  (.D(n_106_642), .CK(n_0), .Q(\mem[61] [2]), .QN());
   DFF_X1 \mem_reg[61][1]  (.D(n_106_641), .CK(n_0), .Q(\mem[61] [1]), .QN());
   DFF_X1 \mem_reg[61][0]  (.D(n_106_640), .CK(n_0), .Q(\mem[61] [0]), .QN());
   DFF_X1 \mem_reg[62][15]  (.D(n_106_639), .CK(n_0), .Q(\mem[62] [15]), .QN());
   DFF_X1 \mem_reg[62][14]  (.D(n_106_638), .CK(n_0), .Q(\mem[62] [14]), .QN());
   DFF_X1 \mem_reg[62][13]  (.D(n_106_637), .CK(n_0), .Q(\mem[62] [13]), .QN());
   DFF_X1 \mem_reg[62][12]  (.D(n_106_636), .CK(n_0), .Q(\mem[62] [12]), .QN());
   DFF_X1 \mem_reg[62][11]  (.D(n_106_635), .CK(n_0), .Q(\mem[62] [11]), .QN());
   DFF_X1 \mem_reg[62][10]  (.D(n_106_634), .CK(n_0), .Q(\mem[62] [10]), .QN());
   DFF_X1 \mem_reg[62][9]  (.D(n_106_633), .CK(n_0), .Q(\mem[62] [9]), .QN());
   DFF_X1 \mem_reg[62][8]  (.D(n_106_632), .CK(n_0), .Q(\mem[62] [8]), .QN());
   DFF_X1 \mem_reg[62][7]  (.D(n_106_631), .CK(n_0), .Q(\mem[62] [7]), .QN());
   DFF_X1 \mem_reg[62][6]  (.D(n_106_630), .CK(n_0), .Q(\mem[62] [6]), .QN());
   DFF_X1 \mem_reg[62][5]  (.D(n_106_629), .CK(n_0), .Q(\mem[62] [5]), .QN());
   DFF_X1 \mem_reg[62][4]  (.D(n_106_628), .CK(n_0), .Q(\mem[62] [4]), .QN());
   DFF_X1 \mem_reg[62][3]  (.D(n_106_627), .CK(n_0), .Q(\mem[62] [3]), .QN());
   DFF_X1 \mem_reg[62][2]  (.D(n_106_626), .CK(n_0), .Q(\mem[62] [2]), .QN());
   DFF_X1 \mem_reg[62][1]  (.D(n_106_625), .CK(n_0), .Q(\mem[62] [1]), .QN());
   DFF_X1 \mem_reg[62][0]  (.D(n_106_624), .CK(n_0), .Q(\mem[62] [0]), .QN());
   DFF_X1 \mem_reg[63][15]  (.D(n_106_623), .CK(n_0), .Q(\mem[63] [15]), .QN());
   DFF_X1 \mem_reg[63][14]  (.D(n_106_622), .CK(n_0), .Q(\mem[63] [14]), .QN());
   DFF_X1 \mem_reg[63][13]  (.D(n_106_621), .CK(n_0), .Q(\mem[63] [13]), .QN());
   DFF_X1 \mem_reg[63][12]  (.D(n_106_620), .CK(n_0), .Q(\mem[63] [12]), .QN());
   DFF_X1 \mem_reg[63][11]  (.D(n_106_619), .CK(n_0), .Q(\mem[63] [11]), .QN());
   DFF_X1 \mem_reg[63][10]  (.D(n_106_618), .CK(n_0), .Q(\mem[63] [10]), .QN());
   DFF_X1 \mem_reg[63][9]  (.D(n_106_617), .CK(n_0), .Q(\mem[63] [9]), .QN());
   DFF_X1 \mem_reg[63][8]  (.D(n_106_616), .CK(n_0), .Q(\mem[63] [8]), .QN());
   DFF_X1 \mem_reg[63][7]  (.D(n_106_615), .CK(n_0), .Q(\mem[63] [7]), .QN());
   DFF_X1 \mem_reg[63][6]  (.D(n_106_614), .CK(n_0), .Q(\mem[63] [6]), .QN());
   DFF_X1 \mem_reg[63][5]  (.D(n_106_613), .CK(n_0), .Q(\mem[63] [5]), .QN());
   DFF_X1 \mem_reg[63][4]  (.D(n_106_612), .CK(n_0), .Q(\mem[63] [4]), .QN());
   DFF_X1 \mem_reg[63][3]  (.D(n_106_611), .CK(n_0), .Q(\mem[63] [3]), .QN());
   DFF_X1 \mem_reg[63][2]  (.D(n_106_610), .CK(n_0), .Q(\mem[63] [2]), .QN());
   DFF_X1 \mem_reg[63][1]  (.D(n_106_609), .CK(n_0), .Q(\mem[63] [1]), .QN());
   DFF_X1 \mem_reg[63][0]  (.D(n_106_608), .CK(n_0), .Q(\mem[63] [0]), .QN());
   DFF_X1 \mem_reg[64][15]  (.D(n_106_607), .CK(n_0), .Q(\mem[64] [15]), .QN());
   DFF_X1 \mem_reg[64][14]  (.D(n_106_606), .CK(n_0), .Q(\mem[64] [14]), .QN());
   DFF_X1 \mem_reg[64][13]  (.D(n_106_605), .CK(n_0), .Q(\mem[64] [13]), .QN());
   DFF_X1 \mem_reg[64][12]  (.D(n_106_604), .CK(n_0), .Q(\mem[64] [12]), .QN());
   DFF_X1 \mem_reg[64][11]  (.D(n_106_603), .CK(n_0), .Q(\mem[64] [11]), .QN());
   DFF_X1 \mem_reg[64][10]  (.D(n_106_602), .CK(n_0), .Q(\mem[64] [10]), .QN());
   DFF_X1 \mem_reg[64][9]  (.D(n_106_601), .CK(n_0), .Q(\mem[64] [9]), .QN());
   DFF_X1 \mem_reg[64][8]  (.D(n_106_600), .CK(n_0), .Q(\mem[64] [8]), .QN());
   DFF_X1 \mem_reg[64][7]  (.D(n_106_599), .CK(n_0), .Q(\mem[64] [7]), .QN());
   DFF_X1 \mem_reg[64][6]  (.D(n_106_598), .CK(n_0), .Q(\mem[64] [6]), .QN());
   DFF_X1 \mem_reg[64][5]  (.D(n_106_597), .CK(n_0), .Q(\mem[64] [5]), .QN());
   DFF_X1 \mem_reg[64][4]  (.D(n_106_596), .CK(n_0), .Q(\mem[64] [4]), .QN());
   DFF_X1 \mem_reg[64][3]  (.D(n_106_595), .CK(n_0), .Q(\mem[64] [3]), .QN());
   DFF_X1 \mem_reg[64][2]  (.D(n_106_594), .CK(n_0), .Q(\mem[64] [2]), .QN());
   DFF_X1 \mem_reg[64][1]  (.D(n_106_593), .CK(n_0), .Q(\mem[64] [1]), .QN());
   DFF_X1 \mem_reg[64][0]  (.D(n_106_592), .CK(n_0), .Q(\mem[64] [0]), .QN());
   DFF_X1 \mem_reg[65][15]  (.D(n_106_591), .CK(n_0), .Q(\mem[65] [15]), .QN());
   DFF_X1 \mem_reg[65][14]  (.D(n_106_590), .CK(n_0), .Q(\mem[65] [14]), .QN());
   DFF_X1 \mem_reg[65][13]  (.D(n_106_589), .CK(n_0), .Q(\mem[65] [13]), .QN());
   DFF_X1 \mem_reg[65][12]  (.D(n_106_588), .CK(n_0), .Q(\mem[65] [12]), .QN());
   DFF_X1 \mem_reg[65][11]  (.D(n_106_587), .CK(n_0), .Q(\mem[65] [11]), .QN());
   DFF_X1 \mem_reg[65][10]  (.D(n_106_586), .CK(n_0), .Q(\mem[65] [10]), .QN());
   DFF_X1 \mem_reg[65][9]  (.D(n_106_585), .CK(n_0), .Q(\mem[65] [9]), .QN());
   DFF_X1 \mem_reg[65][8]  (.D(n_106_584), .CK(n_0), .Q(\mem[65] [8]), .QN());
   DFF_X1 \mem_reg[65][7]  (.D(n_106_583), .CK(n_0), .Q(\mem[65] [7]), .QN());
   DFF_X1 \mem_reg[65][6]  (.D(n_106_582), .CK(n_0), .Q(\mem[65] [6]), .QN());
   DFF_X1 \mem_reg[65][5]  (.D(n_106_581), .CK(n_0), .Q(\mem[65] [5]), .QN());
   DFF_X1 \mem_reg[65][4]  (.D(n_106_580), .CK(n_0), .Q(\mem[65] [4]), .QN());
   DFF_X1 \mem_reg[65][3]  (.D(n_106_579), .CK(n_0), .Q(\mem[65] [3]), .QN());
   DFF_X1 \mem_reg[65][2]  (.D(n_106_578), .CK(n_0), .Q(\mem[65] [2]), .QN());
   DFF_X1 \mem_reg[65][1]  (.D(n_106_577), .CK(n_0), .Q(\mem[65] [1]), .QN());
   DFF_X1 \mem_reg[65][0]  (.D(n_106_576), .CK(n_0), .Q(\mem[65] [0]), .QN());
   DFF_X1 \mem_reg[66][15]  (.D(n_106_575), .CK(n_0), .Q(\mem[66] [15]), .QN());
   DFF_X1 \mem_reg[66][14]  (.D(n_106_574), .CK(n_0), .Q(\mem[66] [14]), .QN());
   DFF_X1 \mem_reg[66][13]  (.D(n_106_573), .CK(n_0), .Q(\mem[66] [13]), .QN());
   DFF_X1 \mem_reg[66][12]  (.D(n_106_572), .CK(n_0), .Q(\mem[66] [12]), .QN());
   DFF_X1 \mem_reg[66][11]  (.D(n_106_571), .CK(n_0), .Q(\mem[66] [11]), .QN());
   DFF_X1 \mem_reg[66][10]  (.D(n_106_570), .CK(n_0), .Q(\mem[66] [10]), .QN());
   DFF_X1 \mem_reg[66][9]  (.D(n_106_569), .CK(n_0), .Q(\mem[66] [9]), .QN());
   DFF_X1 \mem_reg[66][8]  (.D(n_106_568), .CK(n_0), .Q(\mem[66] [8]), .QN());
   DFF_X1 \mem_reg[66][7]  (.D(n_106_567), .CK(n_0), .Q(\mem[66] [7]), .QN());
   DFF_X1 \mem_reg[66][6]  (.D(n_106_566), .CK(n_0), .Q(\mem[66] [6]), .QN());
   DFF_X1 \mem_reg[66][5]  (.D(n_106_565), .CK(n_0), .Q(\mem[66] [5]), .QN());
   DFF_X1 \mem_reg[66][4]  (.D(n_106_564), .CK(n_0), .Q(\mem[66] [4]), .QN());
   DFF_X1 \mem_reg[66][3]  (.D(n_106_563), .CK(n_0), .Q(\mem[66] [3]), .QN());
   DFF_X1 \mem_reg[66][2]  (.D(n_106_562), .CK(n_0), .Q(\mem[66] [2]), .QN());
   DFF_X1 \mem_reg[66][1]  (.D(n_106_561), .CK(n_0), .Q(\mem[66] [1]), .QN());
   DFF_X1 \mem_reg[66][0]  (.D(n_106_560), .CK(n_0), .Q(\mem[66] [0]), .QN());
   DFF_X1 \mem_reg[67][15]  (.D(n_106_559), .CK(n_0), .Q(\mem[67] [15]), .QN());
   DFF_X1 \mem_reg[67][14]  (.D(n_106_558), .CK(n_0), .Q(\mem[67] [14]), .QN());
   DFF_X1 \mem_reg[67][13]  (.D(n_106_557), .CK(n_0), .Q(\mem[67] [13]), .QN());
   DFF_X1 \mem_reg[67][12]  (.D(n_106_556), .CK(n_0), .Q(\mem[67] [12]), .QN());
   DFF_X1 \mem_reg[67][11]  (.D(n_106_555), .CK(n_0), .Q(\mem[67] [11]), .QN());
   DFF_X1 \mem_reg[67][10]  (.D(n_106_554), .CK(n_0), .Q(\mem[67] [10]), .QN());
   DFF_X1 \mem_reg[67][9]  (.D(n_106_553), .CK(n_0), .Q(\mem[67] [9]), .QN());
   DFF_X1 \mem_reg[67][8]  (.D(n_106_552), .CK(n_0), .Q(\mem[67] [8]), .QN());
   DFF_X1 \mem_reg[67][7]  (.D(n_106_551), .CK(n_0), .Q(\mem[67] [7]), .QN());
   DFF_X1 \mem_reg[67][6]  (.D(n_106_550), .CK(n_0), .Q(\mem[67] [6]), .QN());
   DFF_X1 \mem_reg[67][5]  (.D(n_106_549), .CK(n_0), .Q(\mem[67] [5]), .QN());
   DFF_X1 \mem_reg[67][4]  (.D(n_106_548), .CK(n_0), .Q(\mem[67] [4]), .QN());
   DFF_X1 \mem_reg[67][3]  (.D(n_106_547), .CK(n_0), .Q(\mem[67] [3]), .QN());
   DFF_X1 \mem_reg[67][2]  (.D(n_106_546), .CK(n_0), .Q(\mem[67] [2]), .QN());
   DFF_X1 \mem_reg[67][1]  (.D(n_106_545), .CK(n_0), .Q(\mem[67] [1]), .QN());
   DFF_X1 \mem_reg[67][0]  (.D(n_106_544), .CK(n_0), .Q(\mem[67] [0]), .QN());
   DFF_X1 \mem_reg[68][15]  (.D(n_106_543), .CK(n_0), .Q(\mem[68] [15]), .QN());
   DFF_X1 \mem_reg[68][14]  (.D(n_106_542), .CK(n_0), .Q(\mem[68] [14]), .QN());
   DFF_X1 \mem_reg[68][13]  (.D(n_106_541), .CK(n_0), .Q(\mem[68] [13]), .QN());
   DFF_X1 \mem_reg[68][12]  (.D(n_106_540), .CK(n_0), .Q(\mem[68] [12]), .QN());
   DFF_X1 \mem_reg[68][11]  (.D(n_106_539), .CK(n_0), .Q(\mem[68] [11]), .QN());
   DFF_X1 \mem_reg[68][10]  (.D(n_106_538), .CK(n_0), .Q(\mem[68] [10]), .QN());
   DFF_X1 \mem_reg[68][9]  (.D(n_106_537), .CK(n_0), .Q(\mem[68] [9]), .QN());
   DFF_X1 \mem_reg[68][8]  (.D(n_106_536), .CK(n_0), .Q(\mem[68] [8]), .QN());
   DFF_X1 \mem_reg[68][7]  (.D(n_106_535), .CK(n_0), .Q(\mem[68] [7]), .QN());
   DFF_X1 \mem_reg[68][6]  (.D(n_106_534), .CK(n_0), .Q(\mem[68] [6]), .QN());
   DFF_X1 \mem_reg[68][5]  (.D(n_106_533), .CK(n_0), .Q(\mem[68] [5]), .QN());
   DFF_X1 \mem_reg[68][4]  (.D(n_106_532), .CK(n_0), .Q(\mem[68] [4]), .QN());
   DFF_X1 \mem_reg[68][3]  (.D(n_106_531), .CK(n_0), .Q(\mem[68] [3]), .QN());
   DFF_X1 \mem_reg[68][2]  (.D(n_106_530), .CK(n_0), .Q(\mem[68] [2]), .QN());
   DFF_X1 \mem_reg[68][1]  (.D(n_106_529), .CK(n_0), .Q(\mem[68] [1]), .QN());
   DFF_X1 \mem_reg[68][0]  (.D(n_106_528), .CK(n_0), .Q(\mem[68] [0]), .QN());
   DFF_X1 \mem_reg[69][15]  (.D(n_106_527), .CK(n_0), .Q(\mem[69] [15]), .QN());
   DFF_X1 \mem_reg[69][14]  (.D(n_106_526), .CK(n_0), .Q(\mem[69] [14]), .QN());
   DFF_X1 \mem_reg[69][13]  (.D(n_106_525), .CK(n_0), .Q(\mem[69] [13]), .QN());
   DFF_X1 \mem_reg[69][12]  (.D(n_106_524), .CK(n_0), .Q(\mem[69] [12]), .QN());
   DFF_X1 \mem_reg[69][11]  (.D(n_106_523), .CK(n_0), .Q(\mem[69] [11]), .QN());
   DFF_X1 \mem_reg[69][10]  (.D(n_106_522), .CK(n_0), .Q(\mem[69] [10]), .QN());
   DFF_X1 \mem_reg[69][9]  (.D(n_106_521), .CK(n_0), .Q(\mem[69] [9]), .QN());
   DFF_X1 \mem_reg[69][8]  (.D(n_106_520), .CK(n_0), .Q(\mem[69] [8]), .QN());
   DFF_X1 \mem_reg[69][7]  (.D(n_106_519), .CK(n_0), .Q(\mem[69] [7]), .QN());
   DFF_X1 \mem_reg[69][6]  (.D(n_106_518), .CK(n_0), .Q(\mem[69] [6]), .QN());
   DFF_X1 \mem_reg[69][5]  (.D(n_106_517), .CK(n_0), .Q(\mem[69] [5]), .QN());
   DFF_X1 \mem_reg[69][4]  (.D(n_106_516), .CK(n_0), .Q(\mem[69] [4]), .QN());
   DFF_X1 \mem_reg[69][3]  (.D(n_106_515), .CK(n_0), .Q(\mem[69] [3]), .QN());
   DFF_X1 \mem_reg[69][2]  (.D(n_106_514), .CK(n_0), .Q(\mem[69] [2]), .QN());
   DFF_X1 \mem_reg[69][1]  (.D(n_106_513), .CK(n_0), .Q(\mem[69] [1]), .QN());
   DFF_X1 \mem_reg[69][0]  (.D(n_106_512), .CK(n_0), .Q(\mem[69] [0]), .QN());
   DFF_X1 \mem_reg[70][15]  (.D(n_106_511), .CK(n_0), .Q(\mem[70] [15]), .QN());
   DFF_X1 \mem_reg[70][14]  (.D(n_106_510), .CK(n_0), .Q(\mem[70] [14]), .QN());
   DFF_X1 \mem_reg[70][13]  (.D(n_106_509), .CK(n_0), .Q(\mem[70] [13]), .QN());
   DFF_X1 \mem_reg[70][12]  (.D(n_106_508), .CK(n_0), .Q(\mem[70] [12]), .QN());
   DFF_X1 \mem_reg[70][11]  (.D(n_106_507), .CK(n_0), .Q(\mem[70] [11]), .QN());
   DFF_X1 \mem_reg[70][10]  (.D(n_106_506), .CK(n_0), .Q(\mem[70] [10]), .QN());
   DFF_X1 \mem_reg[70][9]  (.D(n_106_505), .CK(n_0), .Q(\mem[70] [9]), .QN());
   DFF_X1 \mem_reg[70][8]  (.D(n_106_504), .CK(n_0), .Q(\mem[70] [8]), .QN());
   DFF_X1 \mem_reg[70][7]  (.D(n_106_503), .CK(n_0), .Q(\mem[70] [7]), .QN());
   DFF_X1 \mem_reg[70][6]  (.D(n_106_502), .CK(n_0), .Q(\mem[70] [6]), .QN());
   DFF_X1 \mem_reg[70][5]  (.D(n_106_501), .CK(n_0), .Q(\mem[70] [5]), .QN());
   DFF_X1 \mem_reg[70][4]  (.D(n_106_500), .CK(n_0), .Q(\mem[70] [4]), .QN());
   DFF_X1 \mem_reg[70][3]  (.D(n_106_499), .CK(n_0), .Q(\mem[70] [3]), .QN());
   DFF_X1 \mem_reg[70][2]  (.D(n_106_498), .CK(n_0), .Q(\mem[70] [2]), .QN());
   DFF_X1 \mem_reg[70][1]  (.D(n_106_497), .CK(n_0), .Q(\mem[70] [1]), .QN());
   DFF_X1 \mem_reg[70][0]  (.D(n_106_496), .CK(n_0), .Q(\mem[70] [0]), .QN());
   DFF_X1 \mem_reg[71][15]  (.D(n_106_495), .CK(n_0), .Q(\mem[71] [15]), .QN());
   DFF_X1 \mem_reg[71][14]  (.D(n_106_494), .CK(n_0), .Q(\mem[71] [14]), .QN());
   DFF_X1 \mem_reg[71][13]  (.D(n_106_493), .CK(n_0), .Q(\mem[71] [13]), .QN());
   DFF_X1 \mem_reg[71][12]  (.D(n_106_492), .CK(n_0), .Q(\mem[71] [12]), .QN());
   DFF_X1 \mem_reg[71][11]  (.D(n_106_491), .CK(n_0), .Q(\mem[71] [11]), .QN());
   DFF_X1 \mem_reg[71][10]  (.D(n_106_490), .CK(n_0), .Q(\mem[71] [10]), .QN());
   DFF_X1 \mem_reg[71][9]  (.D(n_106_489), .CK(n_0), .Q(\mem[71] [9]), .QN());
   DFF_X1 \mem_reg[71][8]  (.D(n_106_488), .CK(n_0), .Q(\mem[71] [8]), .QN());
   DFF_X1 \mem_reg[71][7]  (.D(n_106_487), .CK(n_0), .Q(\mem[71] [7]), .QN());
   DFF_X1 \mem_reg[71][6]  (.D(n_106_486), .CK(n_0), .Q(\mem[71] [6]), .QN());
   DFF_X1 \mem_reg[71][5]  (.D(n_106_485), .CK(n_0), .Q(\mem[71] [5]), .QN());
   DFF_X1 \mem_reg[71][4]  (.D(n_106_484), .CK(n_0), .Q(\mem[71] [4]), .QN());
   DFF_X1 \mem_reg[71][3]  (.D(n_106_483), .CK(n_0), .Q(\mem[71] [3]), .QN());
   DFF_X1 \mem_reg[71][2]  (.D(n_106_482), .CK(n_0), .Q(\mem[71] [2]), .QN());
   DFF_X1 \mem_reg[71][1]  (.D(n_106_481), .CK(n_0), .Q(\mem[71] [1]), .QN());
   DFF_X1 \mem_reg[71][0]  (.D(n_106_480), .CK(n_0), .Q(\mem[71] [0]), .QN());
   DFF_X1 \mem_reg[72][15]  (.D(n_106_479), .CK(n_0), .Q(\mem[72] [15]), .QN());
   DFF_X1 \mem_reg[72][14]  (.D(n_106_478), .CK(n_0), .Q(\mem[72] [14]), .QN());
   DFF_X1 \mem_reg[72][13]  (.D(n_106_477), .CK(n_0), .Q(\mem[72] [13]), .QN());
   DFF_X1 \mem_reg[72][12]  (.D(n_106_476), .CK(n_0), .Q(\mem[72] [12]), .QN());
   DFF_X1 \mem_reg[72][11]  (.D(n_106_475), .CK(n_0), .Q(\mem[72] [11]), .QN());
   DFF_X1 \mem_reg[72][10]  (.D(n_106_474), .CK(n_0), .Q(\mem[72] [10]), .QN());
   DFF_X1 \mem_reg[72][9]  (.D(n_106_473), .CK(n_0), .Q(\mem[72] [9]), .QN());
   DFF_X1 \mem_reg[72][8]  (.D(n_106_472), .CK(n_0), .Q(\mem[72] [8]), .QN());
   DFF_X1 \mem_reg[72][7]  (.D(n_106_471), .CK(n_0), .Q(\mem[72] [7]), .QN());
   DFF_X1 \mem_reg[72][6]  (.D(n_106_470), .CK(n_0), .Q(\mem[72] [6]), .QN());
   DFF_X1 \mem_reg[72][5]  (.D(n_106_469), .CK(n_0), .Q(\mem[72] [5]), .QN());
   DFF_X1 \mem_reg[72][4]  (.D(n_106_468), .CK(n_0), .Q(\mem[72] [4]), .QN());
   DFF_X1 \mem_reg[72][3]  (.D(n_106_467), .CK(n_0), .Q(\mem[72] [3]), .QN());
   DFF_X1 \mem_reg[72][2]  (.D(n_106_466), .CK(n_0), .Q(\mem[72] [2]), .QN());
   DFF_X1 \mem_reg[72][1]  (.D(n_106_465), .CK(n_0), .Q(\mem[72] [1]), .QN());
   DFF_X1 \mem_reg[72][0]  (.D(n_106_464), .CK(n_0), .Q(\mem[72] [0]), .QN());
   DFF_X1 \mem_reg[73][15]  (.D(n_106_463), .CK(n_0), .Q(\mem[73] [15]), .QN());
   DFF_X1 \mem_reg[73][14]  (.D(n_106_462), .CK(n_0), .Q(\mem[73] [14]), .QN());
   DFF_X1 \mem_reg[73][13]  (.D(n_106_461), .CK(n_0), .Q(\mem[73] [13]), .QN());
   DFF_X1 \mem_reg[73][12]  (.D(n_106_460), .CK(n_0), .Q(\mem[73] [12]), .QN());
   DFF_X1 \mem_reg[73][11]  (.D(n_106_459), .CK(n_0), .Q(\mem[73] [11]), .QN());
   DFF_X1 \mem_reg[73][10]  (.D(n_106_458), .CK(n_0), .Q(\mem[73] [10]), .QN());
   DFF_X1 \mem_reg[73][9]  (.D(n_106_457), .CK(n_0), .Q(\mem[73] [9]), .QN());
   DFF_X1 \mem_reg[73][8]  (.D(n_106_456), .CK(n_0), .Q(\mem[73] [8]), .QN());
   DFF_X1 \mem_reg[73][7]  (.D(n_106_455), .CK(n_0), .Q(\mem[73] [7]), .QN());
   DFF_X1 \mem_reg[73][6]  (.D(n_106_454), .CK(n_0), .Q(\mem[73] [6]), .QN());
   DFF_X1 \mem_reg[73][5]  (.D(n_106_453), .CK(n_0), .Q(\mem[73] [5]), .QN());
   DFF_X1 \mem_reg[73][4]  (.D(n_106_452), .CK(n_0), .Q(\mem[73] [4]), .QN());
   DFF_X1 \mem_reg[73][3]  (.D(n_106_451), .CK(n_0), .Q(\mem[73] [3]), .QN());
   DFF_X1 \mem_reg[73][2]  (.D(n_106_450), .CK(n_0), .Q(\mem[73] [2]), .QN());
   DFF_X1 \mem_reg[73][1]  (.D(n_106_449), .CK(n_0), .Q(\mem[73] [1]), .QN());
   DFF_X1 \mem_reg[73][0]  (.D(n_106_448), .CK(n_0), .Q(\mem[73] [0]), .QN());
   DFF_X1 \mem_reg[74][15]  (.D(n_106_447), .CK(n_0), .Q(\mem[74] [15]), .QN());
   DFF_X1 \mem_reg[74][14]  (.D(n_106_446), .CK(n_0), .Q(\mem[74] [14]), .QN());
   DFF_X1 \mem_reg[74][13]  (.D(n_106_445), .CK(n_0), .Q(\mem[74] [13]), .QN());
   DFF_X1 \mem_reg[74][12]  (.D(n_106_444), .CK(n_0), .Q(\mem[74] [12]), .QN());
   DFF_X1 \mem_reg[74][11]  (.D(n_106_443), .CK(n_0), .Q(\mem[74] [11]), .QN());
   DFF_X1 \mem_reg[74][10]  (.D(n_106_442), .CK(n_0), .Q(\mem[74] [10]), .QN());
   DFF_X1 \mem_reg[74][9]  (.D(n_106_441), .CK(n_0), .Q(\mem[74] [9]), .QN());
   DFF_X1 \mem_reg[74][8]  (.D(n_106_440), .CK(n_0), .Q(\mem[74] [8]), .QN());
   DFF_X1 \mem_reg[74][7]  (.D(n_106_439), .CK(n_0), .Q(\mem[74] [7]), .QN());
   DFF_X1 \mem_reg[74][6]  (.D(n_106_438), .CK(n_0), .Q(\mem[74] [6]), .QN());
   DFF_X1 \mem_reg[74][5]  (.D(n_106_437), .CK(n_0), .Q(\mem[74] [5]), .QN());
   DFF_X1 \mem_reg[74][4]  (.D(n_106_436), .CK(n_0), .Q(\mem[74] [4]), .QN());
   DFF_X1 \mem_reg[74][3]  (.D(n_106_435), .CK(n_0), .Q(\mem[74] [3]), .QN());
   DFF_X1 \mem_reg[74][2]  (.D(n_106_434), .CK(n_0), .Q(\mem[74] [2]), .QN());
   DFF_X1 \mem_reg[74][1]  (.D(n_106_433), .CK(n_0), .Q(\mem[74] [1]), .QN());
   DFF_X1 \mem_reg[74][0]  (.D(n_106_432), .CK(n_0), .Q(\mem[74] [0]), .QN());
   DFF_X1 \mem_reg[75][15]  (.D(n_106_431), .CK(n_0), .Q(\mem[75] [15]), .QN());
   DFF_X1 \mem_reg[75][14]  (.D(n_106_430), .CK(n_0), .Q(\mem[75] [14]), .QN());
   DFF_X1 \mem_reg[75][13]  (.D(n_106_429), .CK(n_0), .Q(\mem[75] [13]), .QN());
   DFF_X1 \mem_reg[75][12]  (.D(n_106_428), .CK(n_0), .Q(\mem[75] [12]), .QN());
   DFF_X1 \mem_reg[75][11]  (.D(n_106_427), .CK(n_0), .Q(\mem[75] [11]), .QN());
   DFF_X1 \mem_reg[75][10]  (.D(n_106_426), .CK(n_0), .Q(\mem[75] [10]), .QN());
   DFF_X1 \mem_reg[75][9]  (.D(n_106_425), .CK(n_0), .Q(\mem[75] [9]), .QN());
   DFF_X1 \mem_reg[75][8]  (.D(n_106_424), .CK(n_0), .Q(\mem[75] [8]), .QN());
   DFF_X1 \mem_reg[75][7]  (.D(n_106_423), .CK(n_0), .Q(\mem[75] [7]), .QN());
   DFF_X1 \mem_reg[75][6]  (.D(n_106_422), .CK(n_0), .Q(\mem[75] [6]), .QN());
   DFF_X1 \mem_reg[75][5]  (.D(n_106_421), .CK(n_0), .Q(\mem[75] [5]), .QN());
   DFF_X1 \mem_reg[75][4]  (.D(n_106_420), .CK(n_0), .Q(\mem[75] [4]), .QN());
   DFF_X1 \mem_reg[75][3]  (.D(n_106_419), .CK(n_0), .Q(\mem[75] [3]), .QN());
   DFF_X1 \mem_reg[75][2]  (.D(n_106_418), .CK(n_0), .Q(\mem[75] [2]), .QN());
   DFF_X1 \mem_reg[75][1]  (.D(n_106_417), .CK(n_0), .Q(\mem[75] [1]), .QN());
   DFF_X1 \mem_reg[75][0]  (.D(n_106_416), .CK(n_0), .Q(\mem[75] [0]), .QN());
   DFF_X1 \mem_reg[76][15]  (.D(n_106_415), .CK(n_0), .Q(\mem[76] [15]), .QN());
   DFF_X1 \mem_reg[76][14]  (.D(n_106_414), .CK(n_0), .Q(\mem[76] [14]), .QN());
   DFF_X1 \mem_reg[76][13]  (.D(n_106_413), .CK(n_0), .Q(\mem[76] [13]), .QN());
   DFF_X1 \mem_reg[76][12]  (.D(n_106_412), .CK(n_0), .Q(\mem[76] [12]), .QN());
   DFF_X1 \mem_reg[76][11]  (.D(n_106_411), .CK(n_0), .Q(\mem[76] [11]), .QN());
   DFF_X1 \mem_reg[76][10]  (.D(n_106_410), .CK(n_0), .Q(\mem[76] [10]), .QN());
   DFF_X1 \mem_reg[76][9]  (.D(n_106_409), .CK(n_0), .Q(\mem[76] [9]), .QN());
   DFF_X1 \mem_reg[76][8]  (.D(n_106_408), .CK(n_0), .Q(\mem[76] [8]), .QN());
   DFF_X1 \mem_reg[76][7]  (.D(n_106_407), .CK(n_0), .Q(\mem[76] [7]), .QN());
   DFF_X1 \mem_reg[76][6]  (.D(n_106_406), .CK(n_0), .Q(\mem[76] [6]), .QN());
   DFF_X1 \mem_reg[76][5]  (.D(n_106_405), .CK(n_0), .Q(\mem[76] [5]), .QN());
   DFF_X1 \mem_reg[76][4]  (.D(n_106_404), .CK(n_0), .Q(\mem[76] [4]), .QN());
   DFF_X1 \mem_reg[76][3]  (.D(n_106_403), .CK(n_0), .Q(\mem[76] [3]), .QN());
   DFF_X1 \mem_reg[76][2]  (.D(n_106_402), .CK(n_0), .Q(\mem[76] [2]), .QN());
   DFF_X1 \mem_reg[76][1]  (.D(n_106_401), .CK(n_0), .Q(\mem[76] [1]), .QN());
   DFF_X1 \mem_reg[76][0]  (.D(n_106_400), .CK(n_0), .Q(\mem[76] [0]), .QN());
   DFF_X1 \mem_reg[77][15]  (.D(n_106_399), .CK(n_0), .Q(\mem[77] [15]), .QN());
   DFF_X1 \mem_reg[77][14]  (.D(n_106_398), .CK(n_0), .Q(\mem[77] [14]), .QN());
   DFF_X1 \mem_reg[77][13]  (.D(n_106_397), .CK(n_0), .Q(\mem[77] [13]), .QN());
   DFF_X1 \mem_reg[77][12]  (.D(n_106_396), .CK(n_0), .Q(\mem[77] [12]), .QN());
   DFF_X1 \mem_reg[77][11]  (.D(n_106_395), .CK(n_0), .Q(\mem[77] [11]), .QN());
   DFF_X1 \mem_reg[77][10]  (.D(n_106_394), .CK(n_0), .Q(\mem[77] [10]), .QN());
   DFF_X1 \mem_reg[77][9]  (.D(n_106_393), .CK(n_0), .Q(\mem[77] [9]), .QN());
   DFF_X1 \mem_reg[77][8]  (.D(n_106_392), .CK(n_0), .Q(\mem[77] [8]), .QN());
   DFF_X1 \mem_reg[77][7]  (.D(n_106_391), .CK(n_0), .Q(\mem[77] [7]), .QN());
   DFF_X1 \mem_reg[77][6]  (.D(n_106_390), .CK(n_0), .Q(\mem[77] [6]), .QN());
   DFF_X1 \mem_reg[77][5]  (.D(n_106_389), .CK(n_0), .Q(\mem[77] [5]), .QN());
   DFF_X1 \mem_reg[77][4]  (.D(n_106_388), .CK(n_0), .Q(\mem[77] [4]), .QN());
   DFF_X1 \mem_reg[77][3]  (.D(n_106_387), .CK(n_0), .Q(\mem[77] [3]), .QN());
   DFF_X1 \mem_reg[77][2]  (.D(n_106_386), .CK(n_0), .Q(\mem[77] [2]), .QN());
   DFF_X1 \mem_reg[77][1]  (.D(n_106_385), .CK(n_0), .Q(\mem[77] [1]), .QN());
   DFF_X1 \mem_reg[77][0]  (.D(n_106_384), .CK(n_0), .Q(\mem[77] [0]), .QN());
   DFF_X1 \mem_reg[78][15]  (.D(n_106_383), .CK(n_0), .Q(\mem[78] [15]), .QN());
   DFF_X1 \mem_reg[78][14]  (.D(n_106_382), .CK(n_0), .Q(\mem[78] [14]), .QN());
   DFF_X1 \mem_reg[78][13]  (.D(n_106_381), .CK(n_0), .Q(\mem[78] [13]), .QN());
   DFF_X1 \mem_reg[78][12]  (.D(n_106_380), .CK(n_0), .Q(\mem[78] [12]), .QN());
   DFF_X1 \mem_reg[78][11]  (.D(n_106_379), .CK(n_0), .Q(\mem[78] [11]), .QN());
   DFF_X1 \mem_reg[78][10]  (.D(n_106_378), .CK(n_0), .Q(\mem[78] [10]), .QN());
   DFF_X1 \mem_reg[78][9]  (.D(n_106_377), .CK(n_0), .Q(\mem[78] [9]), .QN());
   DFF_X1 \mem_reg[78][8]  (.D(n_106_376), .CK(n_0), .Q(\mem[78] [8]), .QN());
   DFF_X1 \mem_reg[78][7]  (.D(n_106_375), .CK(n_0), .Q(\mem[78] [7]), .QN());
   DFF_X1 \mem_reg[78][6]  (.D(n_106_374), .CK(n_0), .Q(\mem[78] [6]), .QN());
   DFF_X1 \mem_reg[78][5]  (.D(n_106_373), .CK(n_0), .Q(\mem[78] [5]), .QN());
   DFF_X1 \mem_reg[78][4]  (.D(n_106_372), .CK(n_0), .Q(\mem[78] [4]), .QN());
   DFF_X1 \mem_reg[78][3]  (.D(n_106_371), .CK(n_0), .Q(\mem[78] [3]), .QN());
   DFF_X1 \mem_reg[78][2]  (.D(n_106_370), .CK(n_0), .Q(\mem[78] [2]), .QN());
   DFF_X1 \mem_reg[78][1]  (.D(n_106_369), .CK(n_0), .Q(\mem[78] [1]), .QN());
   DFF_X1 \mem_reg[78][0]  (.D(n_106_368), .CK(n_0), .Q(\mem[78] [0]), .QN());
   DFF_X1 \mem_reg[79][15]  (.D(n_106_367), .CK(n_0), .Q(\mem[79] [15]), .QN());
   DFF_X1 \mem_reg[79][14]  (.D(n_106_366), .CK(n_0), .Q(\mem[79] [14]), .QN());
   DFF_X1 \mem_reg[79][13]  (.D(n_106_365), .CK(n_0), .Q(\mem[79] [13]), .QN());
   DFF_X1 \mem_reg[79][12]  (.D(n_106_364), .CK(n_0), .Q(\mem[79] [12]), .QN());
   DFF_X1 \mem_reg[79][11]  (.D(n_106_363), .CK(n_0), .Q(\mem[79] [11]), .QN());
   DFF_X1 \mem_reg[79][10]  (.D(n_106_362), .CK(n_0), .Q(\mem[79] [10]), .QN());
   DFF_X1 \mem_reg[79][9]  (.D(n_106_361), .CK(n_0), .Q(\mem[79] [9]), .QN());
   DFF_X1 \mem_reg[79][8]  (.D(n_106_360), .CK(n_0), .Q(\mem[79] [8]), .QN());
   DFF_X1 \mem_reg[79][7]  (.D(n_106_359), .CK(n_0), .Q(\mem[79] [7]), .QN());
   DFF_X1 \mem_reg[79][6]  (.D(n_106_358), .CK(n_0), .Q(\mem[79] [6]), .QN());
   DFF_X1 \mem_reg[79][5]  (.D(n_106_357), .CK(n_0), .Q(\mem[79] [5]), .QN());
   DFF_X1 \mem_reg[79][4]  (.D(n_106_356), .CK(n_0), .Q(\mem[79] [4]), .QN());
   DFF_X1 \mem_reg[79][3]  (.D(n_106_355), .CK(n_0), .Q(\mem[79] [3]), .QN());
   DFF_X1 \mem_reg[79][2]  (.D(n_106_354), .CK(n_0), .Q(\mem[79] [2]), .QN());
   DFF_X1 \mem_reg[79][1]  (.D(n_106_353), .CK(n_0), .Q(\mem[79] [1]), .QN());
   DFF_X1 \mem_reg[79][0]  (.D(n_106_352), .CK(n_0), .Q(\mem[79] [0]), .QN());
   DFF_X1 \mem_reg[80][15]  (.D(n_106_351), .CK(n_0), .Q(\mem[80] [15]), .QN());
   DFF_X1 \mem_reg[80][14]  (.D(n_106_350), .CK(n_0), .Q(\mem[80] [14]), .QN());
   DFF_X1 \mem_reg[80][13]  (.D(n_106_349), .CK(n_0), .Q(\mem[80] [13]), .QN());
   DFF_X1 \mem_reg[80][12]  (.D(n_106_348), .CK(n_0), .Q(\mem[80] [12]), .QN());
   DFF_X1 \mem_reg[80][11]  (.D(n_106_347), .CK(n_0), .Q(\mem[80] [11]), .QN());
   DFF_X1 \mem_reg[80][10]  (.D(n_106_346), .CK(n_0), .Q(\mem[80] [10]), .QN());
   DFF_X1 \mem_reg[80][9]  (.D(n_106_345), .CK(n_0), .Q(\mem[80] [9]), .QN());
   DFF_X1 \mem_reg[80][8]  (.D(n_106_344), .CK(n_0), .Q(\mem[80] [8]), .QN());
   DFF_X1 \mem_reg[80][7]  (.D(n_106_343), .CK(n_0), .Q(\mem[80] [7]), .QN());
   DFF_X1 \mem_reg[80][6]  (.D(n_106_342), .CK(n_0), .Q(\mem[80] [6]), .QN());
   DFF_X1 \mem_reg[80][5]  (.D(n_106_341), .CK(n_0), .Q(\mem[80] [5]), .QN());
   DFF_X1 \mem_reg[80][4]  (.D(n_106_340), .CK(n_0), .Q(\mem[80] [4]), .QN());
   DFF_X1 \mem_reg[80][3]  (.D(n_106_339), .CK(n_0), .Q(\mem[80] [3]), .QN());
   DFF_X1 \mem_reg[80][2]  (.D(n_106_338), .CK(n_0), .Q(\mem[80] [2]), .QN());
   DFF_X1 \mem_reg[80][1]  (.D(n_106_337), .CK(n_0), .Q(\mem[80] [1]), .QN());
   DFF_X1 \mem_reg[80][0]  (.D(n_106_336), .CK(n_0), .Q(\mem[80] [0]), .QN());
   DFF_X1 \mem_reg[81][15]  (.D(n_106_335), .CK(n_0), .Q(\mem[81] [15]), .QN());
   DFF_X1 \mem_reg[81][14]  (.D(n_106_334), .CK(n_0), .Q(\mem[81] [14]), .QN());
   DFF_X1 \mem_reg[81][13]  (.D(n_106_333), .CK(n_0), .Q(\mem[81] [13]), .QN());
   DFF_X1 \mem_reg[81][12]  (.D(n_106_332), .CK(n_0), .Q(\mem[81] [12]), .QN());
   DFF_X1 \mem_reg[81][11]  (.D(n_106_331), .CK(n_0), .Q(\mem[81] [11]), .QN());
   DFF_X1 \mem_reg[81][10]  (.D(n_106_330), .CK(n_0), .Q(\mem[81] [10]), .QN());
   DFF_X1 \mem_reg[81][9]  (.D(n_106_329), .CK(n_0), .Q(\mem[81] [9]), .QN());
   DFF_X1 \mem_reg[81][8]  (.D(n_106_328), .CK(n_0), .Q(\mem[81] [8]), .QN());
   DFF_X1 \mem_reg[81][7]  (.D(n_106_327), .CK(n_0), .Q(\mem[81] [7]), .QN());
   DFF_X1 \mem_reg[81][6]  (.D(n_106_326), .CK(n_0), .Q(\mem[81] [6]), .QN());
   DFF_X1 \mem_reg[81][5]  (.D(n_106_325), .CK(n_0), .Q(\mem[81] [5]), .QN());
   DFF_X1 \mem_reg[81][4]  (.D(n_106_324), .CK(n_0), .Q(\mem[81] [4]), .QN());
   DFF_X1 \mem_reg[81][3]  (.D(n_106_323), .CK(n_0), .Q(\mem[81] [3]), .QN());
   DFF_X1 \mem_reg[81][2]  (.D(n_106_322), .CK(n_0), .Q(\mem[81] [2]), .QN());
   DFF_X1 \mem_reg[81][1]  (.D(n_106_321), .CK(n_0), .Q(\mem[81] [1]), .QN());
   DFF_X1 \mem_reg[81][0]  (.D(n_106_320), .CK(n_0), .Q(\mem[81] [0]), .QN());
   DFF_X1 \mem_reg[82][15]  (.D(n_106_319), .CK(n_0), .Q(\mem[82] [15]), .QN());
   DFF_X1 \mem_reg[82][14]  (.D(n_106_318), .CK(n_0), .Q(\mem[82] [14]), .QN());
   DFF_X1 \mem_reg[82][13]  (.D(n_106_317), .CK(n_0), .Q(\mem[82] [13]), .QN());
   DFF_X1 \mem_reg[82][12]  (.D(n_106_316), .CK(n_0), .Q(\mem[82] [12]), .QN());
   DFF_X1 \mem_reg[82][11]  (.D(n_106_315), .CK(n_0), .Q(\mem[82] [11]), .QN());
   DFF_X1 \mem_reg[82][10]  (.D(n_106_314), .CK(n_0), .Q(\mem[82] [10]), .QN());
   DFF_X1 \mem_reg[82][9]  (.D(n_106_313), .CK(n_0), .Q(\mem[82] [9]), .QN());
   DFF_X1 \mem_reg[82][8]  (.D(n_106_312), .CK(n_0), .Q(\mem[82] [8]), .QN());
   DFF_X1 \mem_reg[82][7]  (.D(n_106_311), .CK(n_0), .Q(\mem[82] [7]), .QN());
   DFF_X1 \mem_reg[82][6]  (.D(n_106_310), .CK(n_0), .Q(\mem[82] [6]), .QN());
   DFF_X1 \mem_reg[82][5]  (.D(n_106_309), .CK(n_0), .Q(\mem[82] [5]), .QN());
   DFF_X1 \mem_reg[82][4]  (.D(n_106_308), .CK(n_0), .Q(\mem[82] [4]), .QN());
   DFF_X1 \mem_reg[82][3]  (.D(n_106_307), .CK(n_0), .Q(\mem[82] [3]), .QN());
   DFF_X1 \mem_reg[82][2]  (.D(n_106_306), .CK(n_0), .Q(\mem[82] [2]), .QN());
   DFF_X1 \mem_reg[82][1]  (.D(n_106_305), .CK(n_0), .Q(\mem[82] [1]), .QN());
   DFF_X1 \mem_reg[82][0]  (.D(n_106_304), .CK(n_0), .Q(\mem[82] [0]), .QN());
   DFF_X1 \mem_reg[83][15]  (.D(n_106_303), .CK(n_0), .Q(\mem[83] [15]), .QN());
   DFF_X1 \mem_reg[83][14]  (.D(n_106_302), .CK(n_0), .Q(\mem[83] [14]), .QN());
   DFF_X1 \mem_reg[83][13]  (.D(n_106_301), .CK(n_0), .Q(\mem[83] [13]), .QN());
   DFF_X1 \mem_reg[83][12]  (.D(n_106_300), .CK(n_0), .Q(\mem[83] [12]), .QN());
   DFF_X1 \mem_reg[83][11]  (.D(n_106_299), .CK(n_0), .Q(\mem[83] [11]), .QN());
   DFF_X1 \mem_reg[83][10]  (.D(n_106_298), .CK(n_0), .Q(\mem[83] [10]), .QN());
   DFF_X1 \mem_reg[83][9]  (.D(n_106_297), .CK(n_0), .Q(\mem[83] [9]), .QN());
   DFF_X1 \mem_reg[83][8]  (.D(n_106_296), .CK(n_0), .Q(\mem[83] [8]), .QN());
   DFF_X1 \mem_reg[83][7]  (.D(n_106_295), .CK(n_0), .Q(\mem[83] [7]), .QN());
   DFF_X1 \mem_reg[83][6]  (.D(n_106_294), .CK(n_0), .Q(\mem[83] [6]), .QN());
   DFF_X1 \mem_reg[83][5]  (.D(n_106_293), .CK(n_0), .Q(\mem[83] [5]), .QN());
   DFF_X1 \mem_reg[83][4]  (.D(n_106_292), .CK(n_0), .Q(\mem[83] [4]), .QN());
   DFF_X1 \mem_reg[83][3]  (.D(n_106_291), .CK(n_0), .Q(\mem[83] [3]), .QN());
   DFF_X1 \mem_reg[83][2]  (.D(n_106_290), .CK(n_0), .Q(\mem[83] [2]), .QN());
   DFF_X1 \mem_reg[83][1]  (.D(n_106_289), .CK(n_0), .Q(\mem[83] [1]), .QN());
   DFF_X1 \mem_reg[83][0]  (.D(n_106_288), .CK(n_0), .Q(\mem[83] [0]), .QN());
   DFF_X1 \mem_reg[84][15]  (.D(n_106_287), .CK(n_0), .Q(\mem[84] [15]), .QN());
   DFF_X1 \mem_reg[84][14]  (.D(n_106_286), .CK(n_0), .Q(\mem[84] [14]), .QN());
   DFF_X1 \mem_reg[84][13]  (.D(n_106_285), .CK(n_0), .Q(\mem[84] [13]), .QN());
   DFF_X1 \mem_reg[84][12]  (.D(n_106_284), .CK(n_0), .Q(\mem[84] [12]), .QN());
   DFF_X1 \mem_reg[84][11]  (.D(n_106_283), .CK(n_0), .Q(\mem[84] [11]), .QN());
   DFF_X1 \mem_reg[84][10]  (.D(n_106_282), .CK(n_0), .Q(\mem[84] [10]), .QN());
   DFF_X1 \mem_reg[84][9]  (.D(n_106_281), .CK(n_0), .Q(\mem[84] [9]), .QN());
   DFF_X1 \mem_reg[84][8]  (.D(n_106_280), .CK(n_0), .Q(\mem[84] [8]), .QN());
   DFF_X1 \mem_reg[84][7]  (.D(n_106_279), .CK(n_0), .Q(\mem[84] [7]), .QN());
   DFF_X1 \mem_reg[84][6]  (.D(n_106_278), .CK(n_0), .Q(\mem[84] [6]), .QN());
   DFF_X1 \mem_reg[84][5]  (.D(n_106_277), .CK(n_0), .Q(\mem[84] [5]), .QN());
   DFF_X1 \mem_reg[84][4]  (.D(n_106_276), .CK(n_0), .Q(\mem[84] [4]), .QN());
   DFF_X1 \mem_reg[84][3]  (.D(n_106_275), .CK(n_0), .Q(\mem[84] [3]), .QN());
   DFF_X1 \mem_reg[84][2]  (.D(n_106_274), .CK(n_0), .Q(\mem[84] [2]), .QN());
   DFF_X1 \mem_reg[84][1]  (.D(n_106_273), .CK(n_0), .Q(\mem[84] [1]), .QN());
   DFF_X1 \mem_reg[84][0]  (.D(n_106_272), .CK(n_0), .Q(\mem[84] [0]), .QN());
   DFF_X1 \mem_reg[85][15]  (.D(n_106_271), .CK(n_0), .Q(\mem[85] [15]), .QN());
   DFF_X1 \mem_reg[85][14]  (.D(n_106_270), .CK(n_0), .Q(\mem[85] [14]), .QN());
   DFF_X1 \mem_reg[85][13]  (.D(n_106_269), .CK(n_0), .Q(\mem[85] [13]), .QN());
   DFF_X1 \mem_reg[85][12]  (.D(n_106_268), .CK(n_0), .Q(\mem[85] [12]), .QN());
   DFF_X1 \mem_reg[85][11]  (.D(n_106_267), .CK(n_0), .Q(\mem[85] [11]), .QN());
   DFF_X1 \mem_reg[85][10]  (.D(n_106_266), .CK(n_0), .Q(\mem[85] [10]), .QN());
   DFF_X1 \mem_reg[85][9]  (.D(n_106_265), .CK(n_0), .Q(\mem[85] [9]), .QN());
   DFF_X1 \mem_reg[85][8]  (.D(n_106_264), .CK(n_0), .Q(\mem[85] [8]), .QN());
   DFF_X1 \mem_reg[85][7]  (.D(n_106_263), .CK(n_0), .Q(\mem[85] [7]), .QN());
   DFF_X1 \mem_reg[85][6]  (.D(n_106_262), .CK(n_0), .Q(\mem[85] [6]), .QN());
   DFF_X1 \mem_reg[85][5]  (.D(n_106_261), .CK(n_0), .Q(\mem[85] [5]), .QN());
   DFF_X1 \mem_reg[85][4]  (.D(n_106_260), .CK(n_0), .Q(\mem[85] [4]), .QN());
   DFF_X1 \mem_reg[85][3]  (.D(n_106_259), .CK(n_0), .Q(\mem[85] [3]), .QN());
   DFF_X1 \mem_reg[85][2]  (.D(n_106_258), .CK(n_0), .Q(\mem[85] [2]), .QN());
   DFF_X1 \mem_reg[85][1]  (.D(n_106_257), .CK(n_0), .Q(\mem[85] [1]), .QN());
   DFF_X1 \mem_reg[85][0]  (.D(n_106_256), .CK(n_0), .Q(\mem[85] [0]), .QN());
   DFF_X1 \mem_reg[86][15]  (.D(n_106_255), .CK(n_0), .Q(\mem[86] [15]), .QN());
   DFF_X1 \mem_reg[86][14]  (.D(n_106_254), .CK(n_0), .Q(\mem[86] [14]), .QN());
   DFF_X1 \mem_reg[86][13]  (.D(n_106_253), .CK(n_0), .Q(\mem[86] [13]), .QN());
   DFF_X1 \mem_reg[86][12]  (.D(n_106_252), .CK(n_0), .Q(\mem[86] [12]), .QN());
   DFF_X1 \mem_reg[86][11]  (.D(n_106_251), .CK(n_0), .Q(\mem[86] [11]), .QN());
   DFF_X1 \mem_reg[86][10]  (.D(n_106_250), .CK(n_0), .Q(\mem[86] [10]), .QN());
   DFF_X1 \mem_reg[86][9]  (.D(n_106_249), .CK(n_0), .Q(\mem[86] [9]), .QN());
   DFF_X1 \mem_reg[86][8]  (.D(n_106_248), .CK(n_0), .Q(\mem[86] [8]), .QN());
   DFF_X1 \mem_reg[86][7]  (.D(n_106_247), .CK(n_0), .Q(\mem[86] [7]), .QN());
   DFF_X1 \mem_reg[86][6]  (.D(n_106_246), .CK(n_0), .Q(\mem[86] [6]), .QN());
   DFF_X1 \mem_reg[86][5]  (.D(n_106_245), .CK(n_0), .Q(\mem[86] [5]), .QN());
   DFF_X1 \mem_reg[86][4]  (.D(n_106_244), .CK(n_0), .Q(\mem[86] [4]), .QN());
   DFF_X1 \mem_reg[86][3]  (.D(n_106_243), .CK(n_0), .Q(\mem[86] [3]), .QN());
   DFF_X1 \mem_reg[86][2]  (.D(n_106_242), .CK(n_0), .Q(\mem[86] [2]), .QN());
   DFF_X1 \mem_reg[86][1]  (.D(n_106_241), .CK(n_0), .Q(\mem[86] [1]), .QN());
   DFF_X1 \mem_reg[86][0]  (.D(n_106_240), .CK(n_0), .Q(\mem[86] [0]), .QN());
   DFF_X1 \mem_reg[87][15]  (.D(n_106_239), .CK(n_0), .Q(\mem[87] [15]), .QN());
   DFF_X1 \mem_reg[87][14]  (.D(n_106_238), .CK(n_0), .Q(\mem[87] [14]), .QN());
   DFF_X1 \mem_reg[87][13]  (.D(n_106_237), .CK(n_0), .Q(\mem[87] [13]), .QN());
   DFF_X1 \mem_reg[87][12]  (.D(n_106_236), .CK(n_0), .Q(\mem[87] [12]), .QN());
   DFF_X1 \mem_reg[87][11]  (.D(n_106_235), .CK(n_0), .Q(\mem[87] [11]), .QN());
   DFF_X1 \mem_reg[87][10]  (.D(n_106_234), .CK(n_0), .Q(\mem[87] [10]), .QN());
   DFF_X1 \mem_reg[87][9]  (.D(n_106_233), .CK(n_0), .Q(\mem[87] [9]), .QN());
   DFF_X1 \mem_reg[87][8]  (.D(n_106_232), .CK(n_0), .Q(\mem[87] [8]), .QN());
   DFF_X1 \mem_reg[87][7]  (.D(n_106_231), .CK(n_0), .Q(\mem[87] [7]), .QN());
   DFF_X1 \mem_reg[87][6]  (.D(n_106_230), .CK(n_0), .Q(\mem[87] [6]), .QN());
   DFF_X1 \mem_reg[87][5]  (.D(n_106_229), .CK(n_0), .Q(\mem[87] [5]), .QN());
   DFF_X1 \mem_reg[87][4]  (.D(n_106_228), .CK(n_0), .Q(\mem[87] [4]), .QN());
   DFF_X1 \mem_reg[87][3]  (.D(n_106_227), .CK(n_0), .Q(\mem[87] [3]), .QN());
   DFF_X1 \mem_reg[87][2]  (.D(n_106_226), .CK(n_0), .Q(\mem[87] [2]), .QN());
   DFF_X1 \mem_reg[87][1]  (.D(n_106_225), .CK(n_0), .Q(\mem[87] [1]), .QN());
   DFF_X1 \mem_reg[87][0]  (.D(n_106_224), .CK(n_0), .Q(\mem[87] [0]), .QN());
   DFF_X1 \mem_reg[88][15]  (.D(n_106_223), .CK(n_0), .Q(\mem[88] [15]), .QN());
   DFF_X1 \mem_reg[88][14]  (.D(n_106_222), .CK(n_0), .Q(\mem[88] [14]), .QN());
   DFF_X1 \mem_reg[88][13]  (.D(n_106_221), .CK(n_0), .Q(\mem[88] [13]), .QN());
   DFF_X1 \mem_reg[88][12]  (.D(n_106_220), .CK(n_0), .Q(\mem[88] [12]), .QN());
   DFF_X1 \mem_reg[88][11]  (.D(n_106_219), .CK(n_0), .Q(\mem[88] [11]), .QN());
   DFF_X1 \mem_reg[88][10]  (.D(n_106_218), .CK(n_0), .Q(\mem[88] [10]), .QN());
   DFF_X1 \mem_reg[88][9]  (.D(n_106_217), .CK(n_0), .Q(\mem[88] [9]), .QN());
   DFF_X1 \mem_reg[88][8]  (.D(n_106_216), .CK(n_0), .Q(\mem[88] [8]), .QN());
   DFF_X1 \mem_reg[88][7]  (.D(n_106_215), .CK(n_0), .Q(\mem[88] [7]), .QN());
   DFF_X1 \mem_reg[88][6]  (.D(n_106_214), .CK(n_0), .Q(\mem[88] [6]), .QN());
   DFF_X1 \mem_reg[88][5]  (.D(n_106_213), .CK(n_0), .Q(\mem[88] [5]), .QN());
   DFF_X1 \mem_reg[88][4]  (.D(n_106_212), .CK(n_0), .Q(\mem[88] [4]), .QN());
   DFF_X1 \mem_reg[88][3]  (.D(n_106_211), .CK(n_0), .Q(\mem[88] [3]), .QN());
   DFF_X1 \mem_reg[88][2]  (.D(n_106_210), .CK(n_0), .Q(\mem[88] [2]), .QN());
   DFF_X1 \mem_reg[88][1]  (.D(n_106_209), .CK(n_0), .Q(\mem[88] [1]), .QN());
   DFF_X1 \mem_reg[88][0]  (.D(n_106_208), .CK(n_0), .Q(\mem[88] [0]), .QN());
   DFF_X1 \mem_reg[89][15]  (.D(n_106_207), .CK(n_0), .Q(\mem[89] [15]), .QN());
   DFF_X1 \mem_reg[89][14]  (.D(n_106_206), .CK(n_0), .Q(\mem[89] [14]), .QN());
   DFF_X1 \mem_reg[89][13]  (.D(n_106_205), .CK(n_0), .Q(\mem[89] [13]), .QN());
   DFF_X1 \mem_reg[89][12]  (.D(n_106_204), .CK(n_0), .Q(\mem[89] [12]), .QN());
   DFF_X1 \mem_reg[89][11]  (.D(n_106_203), .CK(n_0), .Q(\mem[89] [11]), .QN());
   DFF_X1 \mem_reg[89][10]  (.D(n_106_202), .CK(n_0), .Q(\mem[89] [10]), .QN());
   DFF_X1 \mem_reg[89][9]  (.D(n_106_201), .CK(n_0), .Q(\mem[89] [9]), .QN());
   DFF_X1 \mem_reg[89][8]  (.D(n_106_200), .CK(n_0), .Q(\mem[89] [8]), .QN());
   DFF_X1 \mem_reg[89][7]  (.D(n_106_199), .CK(n_0), .Q(\mem[89] [7]), .QN());
   DFF_X1 \mem_reg[89][6]  (.D(n_106_198), .CK(n_0), .Q(\mem[89] [6]), .QN());
   DFF_X1 \mem_reg[89][5]  (.D(n_106_197), .CK(n_0), .Q(\mem[89] [5]), .QN());
   DFF_X1 \mem_reg[89][4]  (.D(n_106_196), .CK(n_0), .Q(\mem[89] [4]), .QN());
   DFF_X1 \mem_reg[89][3]  (.D(n_106_195), .CK(n_0), .Q(\mem[89] [3]), .QN());
   DFF_X1 \mem_reg[89][2]  (.D(n_106_194), .CK(n_0), .Q(\mem[89] [2]), .QN());
   DFF_X1 \mem_reg[89][1]  (.D(n_106_193), .CK(n_0), .Q(\mem[89] [1]), .QN());
   DFF_X1 \mem_reg[89][0]  (.D(n_106_192), .CK(n_0), .Q(\mem[89] [0]), .QN());
   DFF_X1 \mem_reg[90][15]  (.D(n_106_191), .CK(n_0), .Q(\mem[90] [15]), .QN());
   DFF_X1 \mem_reg[90][14]  (.D(n_106_190), .CK(n_0), .Q(\mem[90] [14]), .QN());
   DFF_X1 \mem_reg[90][13]  (.D(n_106_189), .CK(n_0), .Q(\mem[90] [13]), .QN());
   DFF_X1 \mem_reg[90][12]  (.D(n_106_188), .CK(n_0), .Q(\mem[90] [12]), .QN());
   DFF_X1 \mem_reg[90][11]  (.D(n_106_187), .CK(n_0), .Q(\mem[90] [11]), .QN());
   DFF_X1 \mem_reg[90][10]  (.D(n_106_186), .CK(n_0), .Q(\mem[90] [10]), .QN());
   DFF_X1 \mem_reg[90][9]  (.D(n_106_185), .CK(n_0), .Q(\mem[90] [9]), .QN());
   DFF_X1 \mem_reg[90][8]  (.D(n_106_184), .CK(n_0), .Q(\mem[90] [8]), .QN());
   DFF_X1 \mem_reg[90][7]  (.D(n_106_183), .CK(n_0), .Q(\mem[90] [7]), .QN());
   DFF_X1 \mem_reg[90][6]  (.D(n_106_182), .CK(n_0), .Q(\mem[90] [6]), .QN());
   DFF_X1 \mem_reg[90][5]  (.D(n_106_181), .CK(n_0), .Q(\mem[90] [5]), .QN());
   DFF_X1 \mem_reg[90][4]  (.D(n_106_180), .CK(n_0), .Q(\mem[90] [4]), .QN());
   DFF_X1 \mem_reg[90][3]  (.D(n_106_179), .CK(n_0), .Q(\mem[90] [3]), .QN());
   DFF_X1 \mem_reg[90][2]  (.D(n_106_178), .CK(n_0), .Q(\mem[90] [2]), .QN());
   DFF_X1 \mem_reg[90][1]  (.D(n_106_177), .CK(n_0), .Q(\mem[90] [1]), .QN());
   DFF_X1 \mem_reg[90][0]  (.D(n_106_176), .CK(n_0), .Q(\mem[90] [0]), .QN());
   DFF_X1 \mem_reg[91][15]  (.D(n_106_175), .CK(n_0), .Q(\mem[91] [15]), .QN());
   DFF_X1 \mem_reg[91][14]  (.D(n_106_174), .CK(n_0), .Q(\mem[91] [14]), .QN());
   DFF_X1 \mem_reg[91][13]  (.D(n_106_173), .CK(n_0), .Q(\mem[91] [13]), .QN());
   DFF_X1 \mem_reg[91][12]  (.D(n_106_172), .CK(n_0), .Q(\mem[91] [12]), .QN());
   DFF_X1 \mem_reg[91][11]  (.D(n_106_171), .CK(n_0), .Q(\mem[91] [11]), .QN());
   DFF_X1 \mem_reg[91][10]  (.D(n_106_170), .CK(n_0), .Q(\mem[91] [10]), .QN());
   DFF_X1 \mem_reg[91][9]  (.D(n_106_169), .CK(n_0), .Q(\mem[91] [9]), .QN());
   DFF_X1 \mem_reg[91][8]  (.D(n_106_168), .CK(n_0), .Q(\mem[91] [8]), .QN());
   DFF_X1 \mem_reg[91][7]  (.D(n_106_167), .CK(n_0), .Q(\mem[91] [7]), .QN());
   DFF_X1 \mem_reg[91][6]  (.D(n_106_166), .CK(n_0), .Q(\mem[91] [6]), .QN());
   DFF_X1 \mem_reg[91][5]  (.D(n_106_165), .CK(n_0), .Q(\mem[91] [5]), .QN());
   DFF_X1 \mem_reg[91][4]  (.D(n_106_164), .CK(n_0), .Q(\mem[91] [4]), .QN());
   DFF_X1 \mem_reg[91][3]  (.D(n_106_163), .CK(n_0), .Q(\mem[91] [3]), .QN());
   DFF_X1 \mem_reg[91][2]  (.D(n_106_162), .CK(n_0), .Q(\mem[91] [2]), .QN());
   DFF_X1 \mem_reg[91][1]  (.D(n_106_161), .CK(n_0), .Q(\mem[91] [1]), .QN());
   DFF_X1 \mem_reg[91][0]  (.D(n_106_160), .CK(n_0), .Q(\mem[91] [0]), .QN());
   DFF_X1 \mem_reg[92][15]  (.D(n_106_159), .CK(n_0), .Q(\mem[92] [15]), .QN());
   DFF_X1 \mem_reg[92][14]  (.D(n_106_158), .CK(n_0), .Q(\mem[92] [14]), .QN());
   DFF_X1 \mem_reg[92][13]  (.D(n_106_157), .CK(n_0), .Q(\mem[92] [13]), .QN());
   DFF_X1 \mem_reg[92][12]  (.D(n_106_156), .CK(n_0), .Q(\mem[92] [12]), .QN());
   DFF_X1 \mem_reg[92][11]  (.D(n_106_155), .CK(n_0), .Q(\mem[92] [11]), .QN());
   DFF_X1 \mem_reg[92][10]  (.D(n_106_154), .CK(n_0), .Q(\mem[92] [10]), .QN());
   DFF_X1 \mem_reg[92][9]  (.D(n_106_153), .CK(n_0), .Q(\mem[92] [9]), .QN());
   DFF_X1 \mem_reg[92][8]  (.D(n_106_152), .CK(n_0), .Q(\mem[92] [8]), .QN());
   DFF_X1 \mem_reg[92][7]  (.D(n_106_151), .CK(n_0), .Q(\mem[92] [7]), .QN());
   DFF_X1 \mem_reg[92][6]  (.D(n_106_150), .CK(n_0), .Q(\mem[92] [6]), .QN());
   DFF_X1 \mem_reg[92][5]  (.D(n_106_149), .CK(n_0), .Q(\mem[92] [5]), .QN());
   DFF_X1 \mem_reg[92][4]  (.D(n_106_148), .CK(n_0), .Q(\mem[92] [4]), .QN());
   DFF_X1 \mem_reg[92][3]  (.D(n_106_147), .CK(n_0), .Q(\mem[92] [3]), .QN());
   DFF_X1 \mem_reg[92][2]  (.D(n_106_146), .CK(n_0), .Q(\mem[92] [2]), .QN());
   DFF_X1 \mem_reg[92][1]  (.D(n_106_145), .CK(n_0), .Q(\mem[92] [1]), .QN());
   DFF_X1 \mem_reg[92][0]  (.D(n_106_144), .CK(n_0), .Q(\mem[92] [0]), .QN());
   DFF_X1 \mem_reg[93][15]  (.D(n_106_143), .CK(n_0), .Q(\mem[93] [15]), .QN());
   DFF_X1 \mem_reg[93][14]  (.D(n_106_142), .CK(n_0), .Q(\mem[93] [14]), .QN());
   DFF_X1 \mem_reg[93][13]  (.D(n_106_141), .CK(n_0), .Q(\mem[93] [13]), .QN());
   DFF_X1 \mem_reg[93][12]  (.D(n_106_140), .CK(n_0), .Q(\mem[93] [12]), .QN());
   DFF_X1 \mem_reg[93][11]  (.D(n_106_139), .CK(n_0), .Q(\mem[93] [11]), .QN());
   DFF_X1 \mem_reg[93][10]  (.D(n_106_138), .CK(n_0), .Q(\mem[93] [10]), .QN());
   DFF_X1 \mem_reg[93][9]  (.D(n_106_137), .CK(n_0), .Q(\mem[93] [9]), .QN());
   DFF_X1 \mem_reg[93][8]  (.D(n_106_136), .CK(n_0), .Q(\mem[93] [8]), .QN());
   DFF_X1 \mem_reg[93][7]  (.D(n_106_135), .CK(n_0), .Q(\mem[93] [7]), .QN());
   DFF_X1 \mem_reg[93][6]  (.D(n_106_134), .CK(n_0), .Q(\mem[93] [6]), .QN());
   DFF_X1 \mem_reg[93][5]  (.D(n_106_133), .CK(n_0), .Q(\mem[93] [5]), .QN());
   DFF_X1 \mem_reg[93][4]  (.D(n_106_132), .CK(n_0), .Q(\mem[93] [4]), .QN());
   DFF_X1 \mem_reg[93][3]  (.D(n_106_131), .CK(n_0), .Q(\mem[93] [3]), .QN());
   DFF_X1 \mem_reg[93][2]  (.D(n_106_130), .CK(n_0), .Q(\mem[93] [2]), .QN());
   DFF_X1 \mem_reg[93][1]  (.D(n_106_129), .CK(n_0), .Q(\mem[93] [1]), .QN());
   DFF_X1 \mem_reg[93][0]  (.D(n_106_128), .CK(n_0), .Q(\mem[93] [0]), .QN());
   DFF_X1 \mem_reg[94][15]  (.D(n_106_127), .CK(n_0), .Q(\mem[94] [15]), .QN());
   DFF_X1 \mem_reg[94][14]  (.D(n_106_126), .CK(n_0), .Q(\mem[94] [14]), .QN());
   DFF_X1 \mem_reg[94][13]  (.D(n_106_125), .CK(n_0), .Q(\mem[94] [13]), .QN());
   DFF_X1 \mem_reg[94][12]  (.D(n_106_124), .CK(n_0), .Q(\mem[94] [12]), .QN());
   DFF_X1 \mem_reg[94][11]  (.D(n_106_123), .CK(n_0), .Q(\mem[94] [11]), .QN());
   DFF_X1 \mem_reg[94][10]  (.D(n_106_122), .CK(n_0), .Q(\mem[94] [10]), .QN());
   DFF_X1 \mem_reg[94][9]  (.D(n_106_121), .CK(n_0), .Q(\mem[94] [9]), .QN());
   DFF_X1 \mem_reg[94][8]  (.D(n_106_120), .CK(n_0), .Q(\mem[94] [8]), .QN());
   DFF_X1 \mem_reg[94][7]  (.D(n_106_119), .CK(n_0), .Q(\mem[94] [7]), .QN());
   DFF_X1 \mem_reg[94][6]  (.D(n_106_118), .CK(n_0), .Q(\mem[94] [6]), .QN());
   DFF_X1 \mem_reg[94][5]  (.D(n_106_117), .CK(n_0), .Q(\mem[94] [5]), .QN());
   DFF_X1 \mem_reg[94][4]  (.D(n_106_116), .CK(n_0), .Q(\mem[94] [4]), .QN());
   DFF_X1 \mem_reg[94][3]  (.D(n_106_115), .CK(n_0), .Q(\mem[94] [3]), .QN());
   DFF_X1 \mem_reg[94][2]  (.D(n_106_114), .CK(n_0), .Q(\mem[94] [2]), .QN());
   DFF_X1 \mem_reg[94][1]  (.D(n_106_113), .CK(n_0), .Q(\mem[94] [1]), .QN());
   DFF_X1 \mem_reg[94][0]  (.D(n_106_112), .CK(n_0), .Q(\mem[94] [0]), .QN());
   DFF_X1 \mem_reg[95][15]  (.D(n_106_111), .CK(n_0), .Q(\mem[95] [15]), .QN());
   DFF_X1 \mem_reg[95][14]  (.D(n_106_110), .CK(n_0), .Q(\mem[95] [14]), .QN());
   DFF_X1 \mem_reg[95][13]  (.D(n_106_109), .CK(n_0), .Q(\mem[95] [13]), .QN());
   DFF_X1 \mem_reg[95][12]  (.D(n_106_108), .CK(n_0), .Q(\mem[95] [12]), .QN());
   DFF_X1 \mem_reg[95][11]  (.D(n_106_107), .CK(n_0), .Q(\mem[95] [11]), .QN());
   DFF_X1 \mem_reg[95][10]  (.D(n_106_106), .CK(n_0), .Q(\mem[95] [10]), .QN());
   DFF_X1 \mem_reg[95][9]  (.D(n_106_105), .CK(n_0), .Q(\mem[95] [9]), .QN());
   DFF_X1 \mem_reg[95][8]  (.D(n_106_104), .CK(n_0), .Q(\mem[95] [8]), .QN());
   DFF_X1 \mem_reg[95][7]  (.D(n_106_103), .CK(n_0), .Q(\mem[95] [7]), .QN());
   DFF_X1 \mem_reg[95][6]  (.D(n_106_102), .CK(n_0), .Q(\mem[95] [6]), .QN());
   DFF_X1 \mem_reg[95][5]  (.D(n_106_101), .CK(n_0), .Q(\mem[95] [5]), .QN());
   DFF_X1 \mem_reg[95][4]  (.D(n_106_100), .CK(n_0), .Q(\mem[95] [4]), .QN());
   DFF_X1 \mem_reg[95][3]  (.D(n_106_99), .CK(n_0), .Q(\mem[95] [3]), .QN());
   DFF_X1 \mem_reg[95][2]  (.D(n_106_98), .CK(n_0), .Q(\mem[95] [2]), .QN());
   DFF_X1 \mem_reg[95][1]  (.D(n_106_97), .CK(n_0), .Q(\mem[95] [1]), .QN());
   DFF_X1 \mem_reg[95][0]  (.D(n_106_96), .CK(n_0), .Q(\mem[95] [0]), .QN());
   DFF_X1 \mem_reg[96][15]  (.D(n_106_95), .CK(n_0), .Q(\mem[96] [15]), .QN());
   DFF_X1 \mem_reg[96][14]  (.D(n_106_94), .CK(n_0), .Q(\mem[96] [14]), .QN());
   DFF_X1 \mem_reg[96][13]  (.D(n_106_93), .CK(n_0), .Q(\mem[96] [13]), .QN());
   DFF_X1 \mem_reg[96][12]  (.D(n_106_92), .CK(n_0), .Q(\mem[96] [12]), .QN());
   DFF_X1 \mem_reg[96][11]  (.D(n_106_91), .CK(n_0), .Q(\mem[96] [11]), .QN());
   DFF_X1 \mem_reg[96][10]  (.D(n_106_90), .CK(n_0), .Q(\mem[96] [10]), .QN());
   DFF_X1 \mem_reg[96][9]  (.D(n_106_89), .CK(n_0), .Q(\mem[96] [9]), .QN());
   DFF_X1 \mem_reg[96][8]  (.D(n_106_88), .CK(n_0), .Q(\mem[96] [8]), .QN());
   DFF_X1 \mem_reg[96][7]  (.D(n_106_87), .CK(n_0), .Q(\mem[96] [7]), .QN());
   DFF_X1 \mem_reg[96][6]  (.D(n_106_86), .CK(n_0), .Q(\mem[96] [6]), .QN());
   DFF_X1 \mem_reg[96][5]  (.D(n_106_85), .CK(n_0), .Q(\mem[96] [5]), .QN());
   DFF_X1 \mem_reg[96][4]  (.D(n_106_84), .CK(n_0), .Q(\mem[96] [4]), .QN());
   DFF_X1 \mem_reg[96][3]  (.D(n_106_83), .CK(n_0), .Q(\mem[96] [3]), .QN());
   DFF_X1 \mem_reg[96][2]  (.D(n_106_82), .CK(n_0), .Q(\mem[96] [2]), .QN());
   DFF_X1 \mem_reg[96][1]  (.D(n_106_81), .CK(n_0), .Q(\mem[96] [1]), .QN());
   DFF_X1 \mem_reg[96][0]  (.D(n_106_80), .CK(n_0), .Q(\mem[96] [0]), .QN());
   DFF_X1 \mem_reg[97][15]  (.D(n_106_79), .CK(n_0), .Q(\mem[97] [15]), .QN());
   DFF_X1 \mem_reg[97][14]  (.D(n_106_78), .CK(n_0), .Q(\mem[97] [14]), .QN());
   DFF_X1 \mem_reg[97][13]  (.D(n_106_77), .CK(n_0), .Q(\mem[97] [13]), .QN());
   DFF_X1 \mem_reg[97][12]  (.D(n_106_76), .CK(n_0), .Q(\mem[97] [12]), .QN());
   DFF_X1 \mem_reg[97][11]  (.D(n_106_75), .CK(n_0), .Q(\mem[97] [11]), .QN());
   DFF_X1 \mem_reg[97][10]  (.D(n_106_74), .CK(n_0), .Q(\mem[97] [10]), .QN());
   DFF_X1 \mem_reg[97][9]  (.D(n_106_73), .CK(n_0), .Q(\mem[97] [9]), .QN());
   DFF_X1 \mem_reg[97][8]  (.D(n_106_72), .CK(n_0), .Q(\mem[97] [8]), .QN());
   DFF_X1 \mem_reg[97][7]  (.D(n_106_71), .CK(n_0), .Q(\mem[97] [7]), .QN());
   DFF_X1 \mem_reg[97][6]  (.D(n_106_70), .CK(n_0), .Q(\mem[97] [6]), .QN());
   DFF_X1 \mem_reg[97][5]  (.D(n_106_69), .CK(n_0), .Q(\mem[97] [5]), .QN());
   DFF_X1 \mem_reg[97][4]  (.D(n_106_68), .CK(n_0), .Q(\mem[97] [4]), .QN());
   DFF_X1 \mem_reg[97][3]  (.D(n_106_67), .CK(n_0), .Q(\mem[97] [3]), .QN());
   DFF_X1 \mem_reg[97][2]  (.D(n_106_66), .CK(n_0), .Q(\mem[97] [2]), .QN());
   DFF_X1 \mem_reg[97][1]  (.D(n_106_65), .CK(n_0), .Q(\mem[97] [1]), .QN());
   DFF_X1 \mem_reg[97][0]  (.D(n_106_64), .CK(n_0), .Q(\mem[97] [0]), .QN());
   DFF_X1 \mem_reg[98][15]  (.D(n_106_63), .CK(n_0), .Q(\mem[98] [15]), .QN());
   DFF_X1 \mem_reg[98][14]  (.D(n_106_62), .CK(n_0), .Q(\mem[98] [14]), .QN());
   DFF_X1 \mem_reg[98][13]  (.D(n_106_61), .CK(n_0), .Q(\mem[98] [13]), .QN());
   DFF_X1 \mem_reg[98][12]  (.D(n_106_60), .CK(n_0), .Q(\mem[98] [12]), .QN());
   DFF_X1 \mem_reg[98][11]  (.D(n_106_59), .CK(n_0), .Q(\mem[98] [11]), .QN());
   DFF_X1 \mem_reg[98][10]  (.D(n_106_58), .CK(n_0), .Q(\mem[98] [10]), .QN());
   DFF_X1 \mem_reg[98][9]  (.D(n_106_57), .CK(n_0), .Q(\mem[98] [9]), .QN());
   DFF_X1 \mem_reg[98][8]  (.D(n_106_56), .CK(n_0), .Q(\mem[98] [8]), .QN());
   DFF_X1 \mem_reg[98][7]  (.D(n_106_55), .CK(n_0), .Q(\mem[98] [7]), .QN());
   DFF_X1 \mem_reg[98][6]  (.D(n_106_54), .CK(n_0), .Q(\mem[98] [6]), .QN());
   DFF_X1 \mem_reg[98][5]  (.D(n_106_53), .CK(n_0), .Q(\mem[98] [5]), .QN());
   DFF_X1 \mem_reg[98][4]  (.D(n_106_52), .CK(n_0), .Q(\mem[98] [4]), .QN());
   DFF_X1 \mem_reg[98][3]  (.D(n_106_51), .CK(n_0), .Q(\mem[98] [3]), .QN());
   DFF_X1 \mem_reg[98][2]  (.D(n_106_50), .CK(n_0), .Q(\mem[98] [2]), .QN());
   DFF_X1 \mem_reg[98][1]  (.D(n_106_49), .CK(n_0), .Q(\mem[98] [1]), .QN());
   DFF_X1 \mem_reg[98][0]  (.D(n_106_48), .CK(n_0), .Q(\mem[98] [0]), .QN());
   DFF_X1 \mem_reg[99][15]  (.D(n_106_47), .CK(n_0), .Q(\mem[99] [15]), .QN());
   DFF_X1 \mem_reg[99][14]  (.D(n_106_46), .CK(n_0), .Q(\mem[99] [14]), .QN());
   DFF_X1 \mem_reg[99][13]  (.D(n_106_45), .CK(n_0), .Q(\mem[99] [13]), .QN());
   DFF_X1 \mem_reg[99][12]  (.D(n_106_44), .CK(n_0), .Q(\mem[99] [12]), .QN());
   DFF_X1 \mem_reg[99][11]  (.D(n_106_43), .CK(n_0), .Q(\mem[99] [11]), .QN());
   DFF_X1 \mem_reg[99][10]  (.D(n_106_42), .CK(n_0), .Q(\mem[99] [10]), .QN());
   DFF_X1 \mem_reg[99][9]  (.D(n_106_41), .CK(n_0), .Q(\mem[99] [9]), .QN());
   DFF_X1 \mem_reg[99][8]  (.D(n_106_40), .CK(n_0), .Q(\mem[99] [8]), .QN());
   DFF_X1 \mem_reg[99][7]  (.D(n_106_39), .CK(n_0), .Q(\mem[99] [7]), .QN());
   DFF_X1 \mem_reg[99][6]  (.D(n_106_38), .CK(n_0), .Q(\mem[99] [6]), .QN());
   DFF_X1 \mem_reg[99][5]  (.D(n_106_37), .CK(n_0), .Q(\mem[99] [5]), .QN());
   DFF_X1 \mem_reg[99][4]  (.D(n_106_36), .CK(n_0), .Q(\mem[99] [4]), .QN());
   DFF_X1 \mem_reg[99][3]  (.D(n_106_35), .CK(n_0), .Q(\mem[99] [3]), .QN());
   DFF_X1 \mem_reg[99][2]  (.D(n_106_34), .CK(n_0), .Q(\mem[99] [2]), .QN());
   DFF_X1 \mem_reg[99][1]  (.D(n_106_33), .CK(n_0), .Q(\mem[99] [1]), .QN());
   DFF_X1 \mem_reg[99][0]  (.D(n_106_32), .CK(n_0), .Q(\mem[99] [0]), .QN());
   DFF_X1 \mem_reg[100][15]  (.D(n_106_31), .CK(n_0), .Q(\mem[100] [15]), .QN());
   DFF_X1 \mem_reg[100][14]  (.D(n_106_30), .CK(n_0), .Q(\mem[100] [14]), .QN());
   DFF_X1 \mem_reg[100][13]  (.D(n_106_29), .CK(n_0), .Q(\mem[100] [13]), .QN());
   DFF_X1 \mem_reg[100][12]  (.D(n_106_28), .CK(n_0), .Q(\mem[100] [12]), .QN());
   DFF_X1 \mem_reg[100][11]  (.D(n_106_27), .CK(n_0), .Q(\mem[100] [11]), .QN());
   DFF_X1 \mem_reg[100][10]  (.D(n_106_26), .CK(n_0), .Q(\mem[100] [10]), .QN());
   DFF_X1 \mem_reg[100][9]  (.D(n_106_25), .CK(n_0), .Q(\mem[100] [9]), .QN());
   DFF_X1 \mem_reg[100][8]  (.D(n_106_24), .CK(n_0), .Q(\mem[100] [8]), .QN());
   DFF_X1 \mem_reg[100][7]  (.D(n_106_23), .CK(n_0), .Q(\mem[100] [7]), .QN());
   DFF_X1 \mem_reg[100][6]  (.D(n_106_22), .CK(n_0), .Q(\mem[100] [6]), .QN());
   DFF_X1 \mem_reg[100][5]  (.D(n_106_21), .CK(n_0), .Q(\mem[100] [5]), .QN());
   DFF_X1 \mem_reg[100][4]  (.D(n_106_20), .CK(n_0), .Q(\mem[100] [4]), .QN());
   DFF_X1 \mem_reg[100][3]  (.D(n_106_19), .CK(n_0), .Q(\mem[100] [3]), .QN());
   DFF_X1 \mem_reg[100][2]  (.D(n_106_18), .CK(n_0), .Q(\mem[100] [2]), .QN());
   DFF_X1 \mem_reg[100][1]  (.D(n_106_17), .CK(n_0), .Q(\mem[100] [1]), .QN());
   DFF_X1 \mem_reg[100][0]  (.D(n_106_16), .CK(n_0), .Q(\mem[100] [0]), .QN());
   DFF_X1 \mem_reg[0][15]  (.D(n_106_15), .CK(n_0), .Q(\mem[0] [15]), .QN());
   DFF_X1 \mem_reg[0][14]  (.D(n_106_14), .CK(n_0), .Q(\mem[0] [14]), .QN());
   DFF_X1 \mem_reg[0][13]  (.D(n_106_13), .CK(n_0), .Q(\mem[0] [13]), .QN());
   DFF_X1 \mem_reg[0][12]  (.D(n_106_12), .CK(n_0), .Q(\mem[0] [12]), .QN());
   DFF_X1 \mem_reg[0][11]  (.D(n_106_11), .CK(n_0), .Q(\mem[0] [11]), .QN());
   DFF_X1 \mem_reg[0][10]  (.D(n_106_10), .CK(n_0), .Q(\mem[0] [10]), .QN());
   DFF_X1 \mem_reg[0][9]  (.D(n_106_9), .CK(n_0), .Q(\mem[0] [9]), .QN());
   DFF_X1 \mem_reg[0][8]  (.D(n_106_8), .CK(n_0), .Q(\mem[0] [8]), .QN());
   DFF_X1 \mem_reg[0][7]  (.D(n_106_7), .CK(n_0), .Q(\mem[0] [7]), .QN());
   DFF_X1 \mem_reg[0][6]  (.D(n_106_6), .CK(n_0), .Q(\mem[0] [6]), .QN());
   DFF_X1 \mem_reg[0][5]  (.D(n_106_5), .CK(n_0), .Q(\mem[0] [5]), .QN());
   DFF_X1 \mem_reg[0][4]  (.D(n_106_4), .CK(n_0), .Q(\mem[0] [4]), .QN());
   DFF_X1 \mem_reg[0][3]  (.D(n_106_3), .CK(n_0), .Q(\mem[0] [3]), .QN());
   DFF_X1 \mem_reg[0][2]  (.D(n_106_2), .CK(n_0), .Q(\mem[0] [2]), .QN());
   DFF_X1 \mem_reg[0][1]  (.D(n_106_1), .CK(n_0), .Q(\mem[0] [1]), .QN());
   DFF_X1 \mem_reg[0][0]  (.D(n_106_0), .CK(n_0), .Q(\mem[0] [0]), .QN());
   MUX2_X1 i_106_0_0 (.A(\mem[52] [15]), .B(data[15]), .S(n_53), .Z(n_106_799));
   MUX2_X1 i_106_0_1 (.A(\mem[52] [14]), .B(data[14]), .S(n_53), .Z(n_106_798));
   MUX2_X1 i_106_0_2 (.A(\mem[52] [13]), .B(data[13]), .S(n_53), .Z(n_106_797));
   MUX2_X1 i_106_0_3 (.A(\mem[52] [12]), .B(data[12]), .S(n_53), .Z(n_106_796));
   MUX2_X1 i_106_0_4 (.A(\mem[52] [11]), .B(data[11]), .S(n_53), .Z(n_106_795));
   MUX2_X1 i_106_0_5 (.A(\mem[52] [10]), .B(data[10]), .S(n_53), .Z(n_106_794));
   MUX2_X1 i_106_0_6 (.A(\mem[52] [9]), .B(data[9]), .S(n_53), .Z(n_106_793));
   MUX2_X1 i_106_0_7 (.A(\mem[52] [8]), .B(data[8]), .S(n_53), .Z(n_106_792));
   MUX2_X1 i_106_0_8 (.A(\mem[52] [7]), .B(data[7]), .S(n_53), .Z(n_106_791));
   MUX2_X1 i_106_0_9 (.A(\mem[52] [6]), .B(data[6]), .S(n_53), .Z(n_106_790));
   MUX2_X1 i_106_0_10 (.A(\mem[52] [5]), .B(data[5]), .S(n_53), .Z(n_106_789));
   MUX2_X1 i_106_0_11 (.A(\mem[52] [4]), .B(data[4]), .S(n_53), .Z(n_106_788));
   MUX2_X1 i_106_0_12 (.A(\mem[52] [3]), .B(data[3]), .S(n_53), .Z(n_106_787));
   MUX2_X1 i_106_0_13 (.A(\mem[52] [2]), .B(data[2]), .S(n_53), .Z(n_106_786));
   MUX2_X1 i_106_0_14 (.A(\mem[52] [1]), .B(data[1]), .S(n_53), .Z(n_106_785));
   MUX2_X1 i_106_0_15 (.A(\mem[52] [0]), .B(data[0]), .S(n_53), .Z(n_106_784));
   MUX2_X1 i_106_0_16 (.A(\mem[53] [15]), .B(data[15]), .S(n_54), .Z(n_106_783));
   MUX2_X1 i_106_0_17 (.A(\mem[53] [14]), .B(data[14]), .S(n_54), .Z(n_106_782));
   MUX2_X1 i_106_0_18 (.A(\mem[53] [13]), .B(data[13]), .S(n_54), .Z(n_106_781));
   MUX2_X1 i_106_0_19 (.A(\mem[53] [12]), .B(data[12]), .S(n_54), .Z(n_106_780));
   MUX2_X1 i_106_0_20 (.A(\mem[53] [11]), .B(data[11]), .S(n_54), .Z(n_106_779));
   MUX2_X1 i_106_0_21 (.A(\mem[53] [10]), .B(data[10]), .S(n_54), .Z(n_106_778));
   MUX2_X1 i_106_0_22 (.A(\mem[53] [9]), .B(data[9]), .S(n_54), .Z(n_106_777));
   MUX2_X1 i_106_0_23 (.A(\mem[53] [8]), .B(data[8]), .S(n_54), .Z(n_106_776));
   MUX2_X1 i_106_0_24 (.A(\mem[53] [7]), .B(data[7]), .S(n_54), .Z(n_106_775));
   MUX2_X1 i_106_0_25 (.A(\mem[53] [6]), .B(data[6]), .S(n_54), .Z(n_106_774));
   MUX2_X1 i_106_0_26 (.A(\mem[53] [5]), .B(data[5]), .S(n_54), .Z(n_106_773));
   MUX2_X1 i_106_0_27 (.A(\mem[53] [4]), .B(data[4]), .S(n_54), .Z(n_106_772));
   MUX2_X1 i_106_0_28 (.A(\mem[53] [3]), .B(data[3]), .S(n_54), .Z(n_106_771));
   MUX2_X1 i_106_0_29 (.A(\mem[53] [2]), .B(data[2]), .S(n_54), .Z(n_106_770));
   MUX2_X1 i_106_0_30 (.A(\mem[53] [1]), .B(data[1]), .S(n_54), .Z(n_106_769));
   MUX2_X1 i_106_0_31 (.A(\mem[53] [0]), .B(data[0]), .S(n_54), .Z(n_106_768));
   MUX2_X1 i_106_0_32 (.A(\mem[54] [15]), .B(data[15]), .S(n_55), .Z(n_106_767));
   MUX2_X1 i_106_0_33 (.A(\mem[54] [14]), .B(data[14]), .S(n_55), .Z(n_106_766));
   MUX2_X1 i_106_0_34 (.A(\mem[54] [13]), .B(data[13]), .S(n_55), .Z(n_106_765));
   MUX2_X1 i_106_0_35 (.A(\mem[54] [12]), .B(data[12]), .S(n_55), .Z(n_106_764));
   MUX2_X1 i_106_0_36 (.A(\mem[54] [11]), .B(data[11]), .S(n_55), .Z(n_106_763));
   MUX2_X1 i_106_0_37 (.A(\mem[54] [10]), .B(data[10]), .S(n_55), .Z(n_106_762));
   MUX2_X1 i_106_0_38 (.A(\mem[54] [9]), .B(data[9]), .S(n_55), .Z(n_106_761));
   MUX2_X1 i_106_0_39 (.A(\mem[54] [8]), .B(data[8]), .S(n_55), .Z(n_106_760));
   MUX2_X1 i_106_0_40 (.A(\mem[54] [7]), .B(data[7]), .S(n_55), .Z(n_106_759));
   MUX2_X1 i_106_0_41 (.A(\mem[54] [6]), .B(data[6]), .S(n_55), .Z(n_106_758));
   MUX2_X1 i_106_0_42 (.A(\mem[54] [5]), .B(data[5]), .S(n_55), .Z(n_106_757));
   MUX2_X1 i_106_0_43 (.A(\mem[54] [4]), .B(data[4]), .S(n_55), .Z(n_106_756));
   MUX2_X1 i_106_0_44 (.A(\mem[54] [3]), .B(data[3]), .S(n_55), .Z(n_106_755));
   MUX2_X1 i_106_0_45 (.A(\mem[54] [2]), .B(data[2]), .S(n_55), .Z(n_106_754));
   MUX2_X1 i_106_0_46 (.A(\mem[54] [1]), .B(data[1]), .S(n_55), .Z(n_106_753));
   MUX2_X1 i_106_0_47 (.A(\mem[54] [0]), .B(data[0]), .S(n_55), .Z(n_106_752));
   MUX2_X1 i_106_0_48 (.A(\mem[55] [15]), .B(data[15]), .S(n_56), .Z(n_106_751));
   MUX2_X1 i_106_0_49 (.A(\mem[55] [14]), .B(data[14]), .S(n_56), .Z(n_106_750));
   MUX2_X1 i_106_0_50 (.A(\mem[55] [13]), .B(data[13]), .S(n_56), .Z(n_106_749));
   MUX2_X1 i_106_0_51 (.A(\mem[55] [12]), .B(data[12]), .S(n_56), .Z(n_106_748));
   MUX2_X1 i_106_0_52 (.A(\mem[55] [11]), .B(data[11]), .S(n_56), .Z(n_106_747));
   MUX2_X1 i_106_0_53 (.A(\mem[55] [10]), .B(data[10]), .S(n_56), .Z(n_106_746));
   MUX2_X1 i_106_0_54 (.A(\mem[55] [9]), .B(data[9]), .S(n_56), .Z(n_106_745));
   MUX2_X1 i_106_0_55 (.A(\mem[55] [8]), .B(data[8]), .S(n_56), .Z(n_106_744));
   MUX2_X1 i_106_0_56 (.A(\mem[55] [7]), .B(data[7]), .S(n_56), .Z(n_106_743));
   MUX2_X1 i_106_0_57 (.A(\mem[55] [6]), .B(data[6]), .S(n_56), .Z(n_106_742));
   MUX2_X1 i_106_0_58 (.A(\mem[55] [5]), .B(data[5]), .S(n_56), .Z(n_106_741));
   MUX2_X1 i_106_0_59 (.A(\mem[55] [4]), .B(data[4]), .S(n_56), .Z(n_106_740));
   MUX2_X1 i_106_0_60 (.A(\mem[55] [3]), .B(data[3]), .S(n_56), .Z(n_106_739));
   MUX2_X1 i_106_0_61 (.A(\mem[55] [2]), .B(data[2]), .S(n_56), .Z(n_106_738));
   MUX2_X1 i_106_0_62 (.A(\mem[55] [1]), .B(data[1]), .S(n_56), .Z(n_106_737));
   MUX2_X1 i_106_0_63 (.A(\mem[55] [0]), .B(data[0]), .S(n_56), .Z(n_106_736));
   MUX2_X1 i_106_0_64 (.A(\mem[56] [15]), .B(data[15]), .S(n_57), .Z(n_106_735));
   MUX2_X1 i_106_0_65 (.A(\mem[56] [14]), .B(data[14]), .S(n_57), .Z(n_106_734));
   MUX2_X1 i_106_0_66 (.A(\mem[56] [13]), .B(data[13]), .S(n_57), .Z(n_106_733));
   MUX2_X1 i_106_0_67 (.A(\mem[56] [12]), .B(data[12]), .S(n_57), .Z(n_106_732));
   MUX2_X1 i_106_0_68 (.A(\mem[56] [11]), .B(data[11]), .S(n_57), .Z(n_106_731));
   MUX2_X1 i_106_0_69 (.A(\mem[56] [10]), .B(data[10]), .S(n_57), .Z(n_106_730));
   MUX2_X1 i_106_0_70 (.A(\mem[56] [9]), .B(data[9]), .S(n_57), .Z(n_106_729));
   MUX2_X1 i_106_0_71 (.A(\mem[56] [8]), .B(data[8]), .S(n_57), .Z(n_106_728));
   MUX2_X1 i_106_0_72 (.A(\mem[56] [7]), .B(data[7]), .S(n_57), .Z(n_106_727));
   MUX2_X1 i_106_0_73 (.A(\mem[56] [6]), .B(data[6]), .S(n_57), .Z(n_106_726));
   MUX2_X1 i_106_0_74 (.A(\mem[56] [5]), .B(data[5]), .S(n_57), .Z(n_106_725));
   MUX2_X1 i_106_0_75 (.A(\mem[56] [4]), .B(data[4]), .S(n_57), .Z(n_106_724));
   MUX2_X1 i_106_0_76 (.A(\mem[56] [3]), .B(data[3]), .S(n_57), .Z(n_106_723));
   MUX2_X1 i_106_0_77 (.A(\mem[56] [2]), .B(data[2]), .S(n_57), .Z(n_106_722));
   MUX2_X1 i_106_0_78 (.A(\mem[56] [1]), .B(data[1]), .S(n_57), .Z(n_106_721));
   MUX2_X1 i_106_0_79 (.A(\mem[56] [0]), .B(data[0]), .S(n_57), .Z(n_106_720));
   MUX2_X1 i_106_0_80 (.A(\mem[57] [15]), .B(data[15]), .S(n_58), .Z(n_106_719));
   MUX2_X1 i_106_0_81 (.A(\mem[57] [14]), .B(data[14]), .S(n_58), .Z(n_106_718));
   MUX2_X1 i_106_0_82 (.A(\mem[57] [13]), .B(data[13]), .S(n_58), .Z(n_106_717));
   MUX2_X1 i_106_0_83 (.A(\mem[57] [12]), .B(data[12]), .S(n_58), .Z(n_106_716));
   MUX2_X1 i_106_0_84 (.A(\mem[57] [11]), .B(data[11]), .S(n_58), .Z(n_106_715));
   MUX2_X1 i_106_0_85 (.A(\mem[57] [10]), .B(data[10]), .S(n_58), .Z(n_106_714));
   MUX2_X1 i_106_0_86 (.A(\mem[57] [9]), .B(data[9]), .S(n_58), .Z(n_106_713));
   MUX2_X1 i_106_0_87 (.A(\mem[57] [8]), .B(data[8]), .S(n_58), .Z(n_106_712));
   MUX2_X1 i_106_0_88 (.A(\mem[57] [7]), .B(data[7]), .S(n_58), .Z(n_106_711));
   MUX2_X1 i_106_0_89 (.A(\mem[57] [6]), .B(data[6]), .S(n_58), .Z(n_106_710));
   MUX2_X1 i_106_0_90 (.A(\mem[57] [5]), .B(data[5]), .S(n_58), .Z(n_106_709));
   MUX2_X1 i_106_0_91 (.A(\mem[57] [4]), .B(data[4]), .S(n_58), .Z(n_106_708));
   MUX2_X1 i_106_0_92 (.A(\mem[57] [3]), .B(data[3]), .S(n_58), .Z(n_106_707));
   MUX2_X1 i_106_0_93 (.A(\mem[57] [2]), .B(data[2]), .S(n_58), .Z(n_106_706));
   MUX2_X1 i_106_0_94 (.A(\mem[57] [1]), .B(data[1]), .S(n_58), .Z(n_106_705));
   MUX2_X1 i_106_0_95 (.A(\mem[57] [0]), .B(data[0]), .S(n_58), .Z(n_106_704));
   MUX2_X1 i_106_0_96 (.A(\mem[58] [15]), .B(data[15]), .S(n_59), .Z(n_106_703));
   MUX2_X1 i_106_0_97 (.A(\mem[58] [14]), .B(data[14]), .S(n_59), .Z(n_106_702));
   MUX2_X1 i_106_0_98 (.A(\mem[58] [13]), .B(data[13]), .S(n_59), .Z(n_106_701));
   MUX2_X1 i_106_0_99 (.A(\mem[58] [12]), .B(data[12]), .S(n_59), .Z(n_106_700));
   MUX2_X1 i_106_0_100 (.A(\mem[58] [11]), .B(data[11]), .S(n_59), .Z(n_106_699));
   MUX2_X1 i_106_0_101 (.A(\mem[58] [10]), .B(data[10]), .S(n_59), .Z(n_106_698));
   MUX2_X1 i_106_0_102 (.A(\mem[58] [9]), .B(data[9]), .S(n_59), .Z(n_106_697));
   MUX2_X1 i_106_0_103 (.A(\mem[58] [8]), .B(data[8]), .S(n_59), .Z(n_106_696));
   MUX2_X1 i_106_0_104 (.A(\mem[58] [7]), .B(data[7]), .S(n_59), .Z(n_106_695));
   MUX2_X1 i_106_0_105 (.A(\mem[58] [6]), .B(data[6]), .S(n_59), .Z(n_106_694));
   MUX2_X1 i_106_0_106 (.A(\mem[58] [5]), .B(data[5]), .S(n_59), .Z(n_106_693));
   MUX2_X1 i_106_0_107 (.A(\mem[58] [4]), .B(data[4]), .S(n_59), .Z(n_106_692));
   MUX2_X1 i_106_0_108 (.A(\mem[58] [3]), .B(data[3]), .S(n_59), .Z(n_106_691));
   MUX2_X1 i_106_0_109 (.A(\mem[58] [2]), .B(data[2]), .S(n_59), .Z(n_106_690));
   MUX2_X1 i_106_0_110 (.A(\mem[58] [1]), .B(data[1]), .S(n_59), .Z(n_106_689));
   MUX2_X1 i_106_0_111 (.A(\mem[58] [0]), .B(data[0]), .S(n_59), .Z(n_106_688));
   MUX2_X1 i_106_0_112 (.A(\mem[59] [15]), .B(data[15]), .S(n_60), .Z(n_106_687));
   MUX2_X1 i_106_0_113 (.A(\mem[59] [14]), .B(data[14]), .S(n_60), .Z(n_106_686));
   MUX2_X1 i_106_0_114 (.A(\mem[59] [13]), .B(data[13]), .S(n_60), .Z(n_106_685));
   MUX2_X1 i_106_0_115 (.A(\mem[59] [12]), .B(data[12]), .S(n_60), .Z(n_106_684));
   MUX2_X1 i_106_0_116 (.A(\mem[59] [11]), .B(data[11]), .S(n_60), .Z(n_106_683));
   MUX2_X1 i_106_0_117 (.A(\mem[59] [10]), .B(data[10]), .S(n_60), .Z(n_106_682));
   MUX2_X1 i_106_0_118 (.A(\mem[59] [9]), .B(data[9]), .S(n_60), .Z(n_106_681));
   MUX2_X1 i_106_0_119 (.A(\mem[59] [8]), .B(data[8]), .S(n_60), .Z(n_106_680));
   MUX2_X1 i_106_0_120 (.A(\mem[59] [7]), .B(data[7]), .S(n_60), .Z(n_106_679));
   MUX2_X1 i_106_0_121 (.A(\mem[59] [6]), .B(data[6]), .S(n_60), .Z(n_106_678));
   MUX2_X1 i_106_0_122 (.A(\mem[59] [5]), .B(data[5]), .S(n_60), .Z(n_106_677));
   MUX2_X1 i_106_0_123 (.A(\mem[59] [4]), .B(data[4]), .S(n_60), .Z(n_106_676));
   MUX2_X1 i_106_0_124 (.A(\mem[59] [3]), .B(data[3]), .S(n_60), .Z(n_106_675));
   MUX2_X1 i_106_0_125 (.A(\mem[59] [2]), .B(data[2]), .S(n_60), .Z(n_106_674));
   MUX2_X1 i_106_0_126 (.A(\mem[59] [1]), .B(data[1]), .S(n_60), .Z(n_106_673));
   MUX2_X1 i_106_0_127 (.A(\mem[59] [0]), .B(data[0]), .S(n_60), .Z(n_106_672));
   MUX2_X1 i_106_0_128 (.A(\mem[60] [15]), .B(data[15]), .S(n_61), .Z(n_106_671));
   MUX2_X1 i_106_0_129 (.A(\mem[60] [14]), .B(data[14]), .S(n_61), .Z(n_106_670));
   MUX2_X1 i_106_0_130 (.A(\mem[60] [13]), .B(data[13]), .S(n_61), .Z(n_106_669));
   MUX2_X1 i_106_0_131 (.A(\mem[60] [12]), .B(data[12]), .S(n_61), .Z(n_106_668));
   MUX2_X1 i_106_0_132 (.A(\mem[60] [11]), .B(data[11]), .S(n_61), .Z(n_106_667));
   MUX2_X1 i_106_0_133 (.A(\mem[60] [10]), .B(data[10]), .S(n_61), .Z(n_106_666));
   MUX2_X1 i_106_0_134 (.A(\mem[60] [9]), .B(data[9]), .S(n_61), .Z(n_106_665));
   MUX2_X1 i_106_0_135 (.A(\mem[60] [8]), .B(data[8]), .S(n_61), .Z(n_106_664));
   MUX2_X1 i_106_0_136 (.A(\mem[60] [7]), .B(data[7]), .S(n_61), .Z(n_106_663));
   MUX2_X1 i_106_0_137 (.A(\mem[60] [6]), .B(data[6]), .S(n_61), .Z(n_106_662));
   MUX2_X1 i_106_0_138 (.A(\mem[60] [5]), .B(data[5]), .S(n_61), .Z(n_106_661));
   MUX2_X1 i_106_0_139 (.A(\mem[60] [4]), .B(data[4]), .S(n_61), .Z(n_106_660));
   MUX2_X1 i_106_0_140 (.A(\mem[60] [3]), .B(data[3]), .S(n_61), .Z(n_106_659));
   MUX2_X1 i_106_0_141 (.A(\mem[60] [2]), .B(data[2]), .S(n_61), .Z(n_106_658));
   MUX2_X1 i_106_0_142 (.A(\mem[60] [1]), .B(data[1]), .S(n_61), .Z(n_106_657));
   MUX2_X1 i_106_0_143 (.A(\mem[60] [0]), .B(data[0]), .S(n_61), .Z(n_106_656));
   MUX2_X1 i_106_0_144 (.A(\mem[61] [15]), .B(data[15]), .S(n_62), .Z(n_106_655));
   MUX2_X1 i_106_0_145 (.A(\mem[61] [14]), .B(data[14]), .S(n_62), .Z(n_106_654));
   MUX2_X1 i_106_0_146 (.A(\mem[61] [13]), .B(data[13]), .S(n_62), .Z(n_106_653));
   MUX2_X1 i_106_0_147 (.A(\mem[61] [12]), .B(data[12]), .S(n_62), .Z(n_106_652));
   MUX2_X1 i_106_0_148 (.A(\mem[61] [11]), .B(data[11]), .S(n_62), .Z(n_106_651));
   MUX2_X1 i_106_0_149 (.A(\mem[61] [10]), .B(data[10]), .S(n_62), .Z(n_106_650));
   MUX2_X1 i_106_0_150 (.A(\mem[61] [9]), .B(data[9]), .S(n_62), .Z(n_106_649));
   MUX2_X1 i_106_0_151 (.A(\mem[61] [8]), .B(data[8]), .S(n_62), .Z(n_106_648));
   MUX2_X1 i_106_0_152 (.A(\mem[61] [7]), .B(data[7]), .S(n_62), .Z(n_106_647));
   MUX2_X1 i_106_0_153 (.A(\mem[61] [6]), .B(data[6]), .S(n_62), .Z(n_106_646));
   MUX2_X1 i_106_0_154 (.A(\mem[61] [5]), .B(data[5]), .S(n_62), .Z(n_106_645));
   MUX2_X1 i_106_0_155 (.A(\mem[61] [4]), .B(data[4]), .S(n_62), .Z(n_106_644));
   MUX2_X1 i_106_0_156 (.A(\mem[61] [3]), .B(data[3]), .S(n_62), .Z(n_106_643));
   MUX2_X1 i_106_0_157 (.A(\mem[61] [2]), .B(data[2]), .S(n_62), .Z(n_106_642));
   MUX2_X1 i_106_0_158 (.A(\mem[61] [1]), .B(data[1]), .S(n_62), .Z(n_106_641));
   MUX2_X1 i_106_0_159 (.A(\mem[61] [0]), .B(data[0]), .S(n_62), .Z(n_106_640));
   MUX2_X1 i_106_0_160 (.A(\mem[62] [15]), .B(data[15]), .S(n_63), .Z(n_106_639));
   MUX2_X1 i_106_0_161 (.A(\mem[62] [14]), .B(data[14]), .S(n_63), .Z(n_106_638));
   MUX2_X1 i_106_0_162 (.A(\mem[62] [13]), .B(data[13]), .S(n_63), .Z(n_106_637));
   MUX2_X1 i_106_0_163 (.A(\mem[62] [12]), .B(data[12]), .S(n_63), .Z(n_106_636));
   MUX2_X1 i_106_0_164 (.A(\mem[62] [11]), .B(data[11]), .S(n_63), .Z(n_106_635));
   MUX2_X1 i_106_0_165 (.A(\mem[62] [10]), .B(data[10]), .S(n_63), .Z(n_106_634));
   MUX2_X1 i_106_0_166 (.A(\mem[62] [9]), .B(data[9]), .S(n_63), .Z(n_106_633));
   MUX2_X1 i_106_0_167 (.A(\mem[62] [8]), .B(data[8]), .S(n_63), .Z(n_106_632));
   MUX2_X1 i_106_0_168 (.A(\mem[62] [7]), .B(data[7]), .S(n_63), .Z(n_106_631));
   MUX2_X1 i_106_0_169 (.A(\mem[62] [6]), .B(data[6]), .S(n_63), .Z(n_106_630));
   MUX2_X1 i_106_0_170 (.A(\mem[62] [5]), .B(data[5]), .S(n_63), .Z(n_106_629));
   MUX2_X1 i_106_0_171 (.A(\mem[62] [4]), .B(data[4]), .S(n_63), .Z(n_106_628));
   MUX2_X1 i_106_0_172 (.A(\mem[62] [3]), .B(data[3]), .S(n_63), .Z(n_106_627));
   MUX2_X1 i_106_0_173 (.A(\mem[62] [2]), .B(data[2]), .S(n_63), .Z(n_106_626));
   MUX2_X1 i_106_0_174 (.A(\mem[62] [1]), .B(data[1]), .S(n_63), .Z(n_106_625));
   MUX2_X1 i_106_0_175 (.A(\mem[62] [0]), .B(data[0]), .S(n_63), .Z(n_106_624));
   MUX2_X1 i_106_0_176 (.A(\mem[63] [15]), .B(data[15]), .S(n_64), .Z(n_106_623));
   MUX2_X1 i_106_0_177 (.A(\mem[63] [14]), .B(data[14]), .S(n_64), .Z(n_106_622));
   MUX2_X1 i_106_0_178 (.A(\mem[63] [13]), .B(data[13]), .S(n_64), .Z(n_106_621));
   MUX2_X1 i_106_0_179 (.A(\mem[63] [12]), .B(data[12]), .S(n_64), .Z(n_106_620));
   MUX2_X1 i_106_0_180 (.A(\mem[63] [11]), .B(data[11]), .S(n_64), .Z(n_106_619));
   MUX2_X1 i_106_0_181 (.A(\mem[63] [10]), .B(data[10]), .S(n_64), .Z(n_106_618));
   MUX2_X1 i_106_0_182 (.A(\mem[63] [9]), .B(data[9]), .S(n_64), .Z(n_106_617));
   MUX2_X1 i_106_0_183 (.A(\mem[63] [8]), .B(data[8]), .S(n_64), .Z(n_106_616));
   MUX2_X1 i_106_0_184 (.A(\mem[63] [7]), .B(data[7]), .S(n_64), .Z(n_106_615));
   MUX2_X1 i_106_0_185 (.A(\mem[63] [6]), .B(data[6]), .S(n_64), .Z(n_106_614));
   MUX2_X1 i_106_0_186 (.A(\mem[63] [5]), .B(data[5]), .S(n_64), .Z(n_106_613));
   MUX2_X1 i_106_0_187 (.A(\mem[63] [4]), .B(data[4]), .S(n_64), .Z(n_106_612));
   MUX2_X1 i_106_0_188 (.A(\mem[63] [3]), .B(data[3]), .S(n_64), .Z(n_106_611));
   MUX2_X1 i_106_0_189 (.A(\mem[63] [2]), .B(data[2]), .S(n_64), .Z(n_106_610));
   MUX2_X1 i_106_0_190 (.A(\mem[63] [1]), .B(data[1]), .S(n_64), .Z(n_106_609));
   MUX2_X1 i_106_0_191 (.A(\mem[63] [0]), .B(data[0]), .S(n_64), .Z(n_106_608));
   MUX2_X1 i_106_0_192 (.A(\mem[64] [15]), .B(data[15]), .S(n_65), .Z(n_106_607));
   MUX2_X1 i_106_0_193 (.A(\mem[64] [14]), .B(data[14]), .S(n_65), .Z(n_106_606));
   MUX2_X1 i_106_0_194 (.A(\mem[64] [13]), .B(data[13]), .S(n_65), .Z(n_106_605));
   MUX2_X1 i_106_0_195 (.A(\mem[64] [12]), .B(data[12]), .S(n_65), .Z(n_106_604));
   MUX2_X1 i_106_0_196 (.A(\mem[64] [11]), .B(data[11]), .S(n_65), .Z(n_106_603));
   MUX2_X1 i_106_0_197 (.A(\mem[64] [10]), .B(data[10]), .S(n_65), .Z(n_106_602));
   MUX2_X1 i_106_0_198 (.A(\mem[64] [9]), .B(data[9]), .S(n_65), .Z(n_106_601));
   MUX2_X1 i_106_0_199 (.A(\mem[64] [8]), .B(data[8]), .S(n_65), .Z(n_106_600));
   MUX2_X1 i_106_0_200 (.A(\mem[64] [7]), .B(data[7]), .S(n_65), .Z(n_106_599));
   MUX2_X1 i_106_0_201 (.A(\mem[64] [6]), .B(data[6]), .S(n_65), .Z(n_106_598));
   MUX2_X1 i_106_0_202 (.A(\mem[64] [5]), .B(data[5]), .S(n_65), .Z(n_106_597));
   MUX2_X1 i_106_0_203 (.A(\mem[64] [4]), .B(data[4]), .S(n_65), .Z(n_106_596));
   MUX2_X1 i_106_0_204 (.A(\mem[64] [3]), .B(data[3]), .S(n_65), .Z(n_106_595));
   MUX2_X1 i_106_0_205 (.A(\mem[64] [2]), .B(data[2]), .S(n_65), .Z(n_106_594));
   MUX2_X1 i_106_0_206 (.A(\mem[64] [1]), .B(data[1]), .S(n_65), .Z(n_106_593));
   MUX2_X1 i_106_0_207 (.A(\mem[64] [0]), .B(data[0]), .S(n_65), .Z(n_106_592));
   MUX2_X1 i_106_0_208 (.A(\mem[65] [15]), .B(data[15]), .S(n_66), .Z(n_106_591));
   MUX2_X1 i_106_0_209 (.A(\mem[65] [14]), .B(data[14]), .S(n_66), .Z(n_106_590));
   MUX2_X1 i_106_0_210 (.A(\mem[65] [13]), .B(data[13]), .S(n_66), .Z(n_106_589));
   MUX2_X1 i_106_0_211 (.A(\mem[65] [12]), .B(data[12]), .S(n_66), .Z(n_106_588));
   MUX2_X1 i_106_0_212 (.A(\mem[65] [11]), .B(data[11]), .S(n_66), .Z(n_106_587));
   MUX2_X1 i_106_0_213 (.A(\mem[65] [10]), .B(data[10]), .S(n_66), .Z(n_106_586));
   MUX2_X1 i_106_0_214 (.A(\mem[65] [9]), .B(data[9]), .S(n_66), .Z(n_106_585));
   MUX2_X1 i_106_0_215 (.A(\mem[65] [8]), .B(data[8]), .S(n_66), .Z(n_106_584));
   MUX2_X1 i_106_0_216 (.A(\mem[65] [7]), .B(data[7]), .S(n_66), .Z(n_106_583));
   MUX2_X1 i_106_0_217 (.A(\mem[65] [6]), .B(data[6]), .S(n_66), .Z(n_106_582));
   MUX2_X1 i_106_0_218 (.A(\mem[65] [5]), .B(data[5]), .S(n_66), .Z(n_106_581));
   MUX2_X1 i_106_0_219 (.A(\mem[65] [4]), .B(data[4]), .S(n_66), .Z(n_106_580));
   MUX2_X1 i_106_0_220 (.A(\mem[65] [3]), .B(data[3]), .S(n_66), .Z(n_106_579));
   MUX2_X1 i_106_0_221 (.A(\mem[65] [2]), .B(data[2]), .S(n_66), .Z(n_106_578));
   MUX2_X1 i_106_0_222 (.A(\mem[65] [1]), .B(data[1]), .S(n_66), .Z(n_106_577));
   MUX2_X1 i_106_0_223 (.A(\mem[65] [0]), .B(data[0]), .S(n_66), .Z(n_106_576));
   MUX2_X1 i_106_0_224 (.A(\mem[66] [15]), .B(data[15]), .S(n_67), .Z(n_106_575));
   MUX2_X1 i_106_0_225 (.A(\mem[66] [14]), .B(data[14]), .S(n_67), .Z(n_106_574));
   MUX2_X1 i_106_0_226 (.A(\mem[66] [13]), .B(data[13]), .S(n_67), .Z(n_106_573));
   MUX2_X1 i_106_0_227 (.A(\mem[66] [12]), .B(data[12]), .S(n_67), .Z(n_106_572));
   MUX2_X1 i_106_0_228 (.A(\mem[66] [11]), .B(data[11]), .S(n_67), .Z(n_106_571));
   MUX2_X1 i_106_0_229 (.A(\mem[66] [10]), .B(data[10]), .S(n_67), .Z(n_106_570));
   MUX2_X1 i_106_0_230 (.A(\mem[66] [9]), .B(data[9]), .S(n_67), .Z(n_106_569));
   MUX2_X1 i_106_0_231 (.A(\mem[66] [8]), .B(data[8]), .S(n_67), .Z(n_106_568));
   MUX2_X1 i_106_0_232 (.A(\mem[66] [7]), .B(data[7]), .S(n_67), .Z(n_106_567));
   MUX2_X1 i_106_0_233 (.A(\mem[66] [6]), .B(data[6]), .S(n_67), .Z(n_106_566));
   MUX2_X1 i_106_0_234 (.A(\mem[66] [5]), .B(data[5]), .S(n_67), .Z(n_106_565));
   MUX2_X1 i_106_0_235 (.A(\mem[66] [4]), .B(data[4]), .S(n_67), .Z(n_106_564));
   MUX2_X1 i_106_0_236 (.A(\mem[66] [3]), .B(data[3]), .S(n_67), .Z(n_106_563));
   MUX2_X1 i_106_0_237 (.A(\mem[66] [2]), .B(data[2]), .S(n_67), .Z(n_106_562));
   MUX2_X1 i_106_0_238 (.A(\mem[66] [1]), .B(data[1]), .S(n_67), .Z(n_106_561));
   MUX2_X1 i_106_0_239 (.A(\mem[66] [0]), .B(data[0]), .S(n_67), .Z(n_106_560));
   MUX2_X1 i_106_0_240 (.A(\mem[67] [15]), .B(data[15]), .S(n_68), .Z(n_106_559));
   MUX2_X1 i_106_0_241 (.A(\mem[67] [14]), .B(data[14]), .S(n_68), .Z(n_106_558));
   MUX2_X1 i_106_0_242 (.A(\mem[67] [13]), .B(data[13]), .S(n_68), .Z(n_106_557));
   MUX2_X1 i_106_0_243 (.A(\mem[67] [12]), .B(data[12]), .S(n_68), .Z(n_106_556));
   MUX2_X1 i_106_0_244 (.A(\mem[67] [11]), .B(data[11]), .S(n_68), .Z(n_106_555));
   MUX2_X1 i_106_0_245 (.A(\mem[67] [10]), .B(data[10]), .S(n_68), .Z(n_106_554));
   MUX2_X1 i_106_0_246 (.A(\mem[67] [9]), .B(data[9]), .S(n_68), .Z(n_106_553));
   MUX2_X1 i_106_0_247 (.A(\mem[67] [8]), .B(data[8]), .S(n_68), .Z(n_106_552));
   MUX2_X1 i_106_0_248 (.A(\mem[67] [7]), .B(data[7]), .S(n_68), .Z(n_106_551));
   MUX2_X1 i_106_0_249 (.A(\mem[67] [6]), .B(data[6]), .S(n_68), .Z(n_106_550));
   MUX2_X1 i_106_0_250 (.A(\mem[67] [5]), .B(data[5]), .S(n_68), .Z(n_106_549));
   MUX2_X1 i_106_0_251 (.A(\mem[67] [4]), .B(data[4]), .S(n_68), .Z(n_106_548));
   MUX2_X1 i_106_0_252 (.A(\mem[67] [3]), .B(data[3]), .S(n_68), .Z(n_106_547));
   MUX2_X1 i_106_0_253 (.A(\mem[67] [2]), .B(data[2]), .S(n_68), .Z(n_106_546));
   MUX2_X1 i_106_0_254 (.A(\mem[67] [1]), .B(data[1]), .S(n_68), .Z(n_106_545));
   MUX2_X1 i_106_0_255 (.A(\mem[67] [0]), .B(data[0]), .S(n_68), .Z(n_106_544));
   MUX2_X1 i_106_0_256 (.A(\mem[68] [15]), .B(data[15]), .S(n_69), .Z(n_106_543));
   MUX2_X1 i_106_0_257 (.A(\mem[68] [14]), .B(data[14]), .S(n_69), .Z(n_106_542));
   MUX2_X1 i_106_0_258 (.A(\mem[68] [13]), .B(data[13]), .S(n_69), .Z(n_106_541));
   MUX2_X1 i_106_0_259 (.A(\mem[68] [12]), .B(data[12]), .S(n_69), .Z(n_106_540));
   MUX2_X1 i_106_0_260 (.A(\mem[68] [11]), .B(data[11]), .S(n_69), .Z(n_106_539));
   MUX2_X1 i_106_0_261 (.A(\mem[68] [10]), .B(data[10]), .S(n_69), .Z(n_106_538));
   MUX2_X1 i_106_0_262 (.A(\mem[68] [9]), .B(data[9]), .S(n_69), .Z(n_106_537));
   MUX2_X1 i_106_0_263 (.A(\mem[68] [8]), .B(data[8]), .S(n_69), .Z(n_106_536));
   MUX2_X1 i_106_0_264 (.A(\mem[68] [7]), .B(data[7]), .S(n_69), .Z(n_106_535));
   MUX2_X1 i_106_0_265 (.A(\mem[68] [6]), .B(data[6]), .S(n_69), .Z(n_106_534));
   MUX2_X1 i_106_0_266 (.A(\mem[68] [5]), .B(data[5]), .S(n_69), .Z(n_106_533));
   MUX2_X1 i_106_0_267 (.A(\mem[68] [4]), .B(data[4]), .S(n_69), .Z(n_106_532));
   MUX2_X1 i_106_0_268 (.A(\mem[68] [3]), .B(data[3]), .S(n_69), .Z(n_106_531));
   MUX2_X1 i_106_0_269 (.A(\mem[68] [2]), .B(data[2]), .S(n_69), .Z(n_106_530));
   MUX2_X1 i_106_0_270 (.A(\mem[68] [1]), .B(data[1]), .S(n_69), .Z(n_106_529));
   MUX2_X1 i_106_0_271 (.A(\mem[68] [0]), .B(data[0]), .S(n_69), .Z(n_106_528));
   MUX2_X1 i_106_0_272 (.A(\mem[69] [15]), .B(data[15]), .S(n_70), .Z(n_106_527));
   MUX2_X1 i_106_0_273 (.A(\mem[69] [14]), .B(data[14]), .S(n_70), .Z(n_106_526));
   MUX2_X1 i_106_0_274 (.A(\mem[69] [13]), .B(data[13]), .S(n_70), .Z(n_106_525));
   MUX2_X1 i_106_0_275 (.A(\mem[69] [12]), .B(data[12]), .S(n_70), .Z(n_106_524));
   MUX2_X1 i_106_0_276 (.A(\mem[69] [11]), .B(data[11]), .S(n_70), .Z(n_106_523));
   MUX2_X1 i_106_0_277 (.A(\mem[69] [10]), .B(data[10]), .S(n_70), .Z(n_106_522));
   MUX2_X1 i_106_0_278 (.A(\mem[69] [9]), .B(data[9]), .S(n_70), .Z(n_106_521));
   MUX2_X1 i_106_0_279 (.A(\mem[69] [8]), .B(data[8]), .S(n_70), .Z(n_106_520));
   MUX2_X1 i_106_0_280 (.A(\mem[69] [7]), .B(data[7]), .S(n_70), .Z(n_106_519));
   MUX2_X1 i_106_0_281 (.A(\mem[69] [6]), .B(data[6]), .S(n_70), .Z(n_106_518));
   MUX2_X1 i_106_0_282 (.A(\mem[69] [5]), .B(data[5]), .S(n_70), .Z(n_106_517));
   MUX2_X1 i_106_0_283 (.A(\mem[69] [4]), .B(data[4]), .S(n_70), .Z(n_106_516));
   MUX2_X1 i_106_0_284 (.A(\mem[69] [3]), .B(data[3]), .S(n_70), .Z(n_106_515));
   MUX2_X1 i_106_0_285 (.A(\mem[69] [2]), .B(data[2]), .S(n_70), .Z(n_106_514));
   MUX2_X1 i_106_0_286 (.A(\mem[69] [1]), .B(data[1]), .S(n_70), .Z(n_106_513));
   MUX2_X1 i_106_0_287 (.A(\mem[69] [0]), .B(data[0]), .S(n_70), .Z(n_106_512));
   MUX2_X1 i_106_0_288 (.A(\mem[70] [15]), .B(data[15]), .S(n_71), .Z(n_106_511));
   MUX2_X1 i_106_0_289 (.A(\mem[70] [14]), .B(data[14]), .S(n_71), .Z(n_106_510));
   MUX2_X1 i_106_0_290 (.A(\mem[70] [13]), .B(data[13]), .S(n_71), .Z(n_106_509));
   MUX2_X1 i_106_0_291 (.A(\mem[70] [12]), .B(data[12]), .S(n_71), .Z(n_106_508));
   MUX2_X1 i_106_0_292 (.A(\mem[70] [11]), .B(data[11]), .S(n_71), .Z(n_106_507));
   MUX2_X1 i_106_0_293 (.A(\mem[70] [10]), .B(data[10]), .S(n_71), .Z(n_106_506));
   MUX2_X1 i_106_0_294 (.A(\mem[70] [9]), .B(data[9]), .S(n_71), .Z(n_106_505));
   MUX2_X1 i_106_0_295 (.A(\mem[70] [8]), .B(data[8]), .S(n_71), .Z(n_106_504));
   MUX2_X1 i_106_0_296 (.A(\mem[70] [7]), .B(data[7]), .S(n_71), .Z(n_106_503));
   MUX2_X1 i_106_0_297 (.A(\mem[70] [6]), .B(data[6]), .S(n_71), .Z(n_106_502));
   MUX2_X1 i_106_0_298 (.A(\mem[70] [5]), .B(data[5]), .S(n_71), .Z(n_106_501));
   MUX2_X1 i_106_0_299 (.A(\mem[70] [4]), .B(data[4]), .S(n_71), .Z(n_106_500));
   MUX2_X1 i_106_0_300 (.A(\mem[70] [3]), .B(data[3]), .S(n_71), .Z(n_106_499));
   MUX2_X1 i_106_0_301 (.A(\mem[70] [2]), .B(data[2]), .S(n_71), .Z(n_106_498));
   MUX2_X1 i_106_0_302 (.A(\mem[70] [1]), .B(data[1]), .S(n_71), .Z(n_106_497));
   MUX2_X1 i_106_0_303 (.A(\mem[70] [0]), .B(data[0]), .S(n_71), .Z(n_106_496));
   MUX2_X1 i_106_0_304 (.A(\mem[71] [15]), .B(data[15]), .S(n_72), .Z(n_106_495));
   MUX2_X1 i_106_0_305 (.A(\mem[71] [14]), .B(data[14]), .S(n_72), .Z(n_106_494));
   MUX2_X1 i_106_0_306 (.A(\mem[71] [13]), .B(data[13]), .S(n_72), .Z(n_106_493));
   MUX2_X1 i_106_0_307 (.A(\mem[71] [12]), .B(data[12]), .S(n_72), .Z(n_106_492));
   MUX2_X1 i_106_0_308 (.A(\mem[71] [11]), .B(data[11]), .S(n_72), .Z(n_106_491));
   MUX2_X1 i_106_0_309 (.A(\mem[71] [10]), .B(data[10]), .S(n_72), .Z(n_106_490));
   MUX2_X1 i_106_0_310 (.A(\mem[71] [9]), .B(data[9]), .S(n_72), .Z(n_106_489));
   MUX2_X1 i_106_0_311 (.A(\mem[71] [8]), .B(data[8]), .S(n_72), .Z(n_106_488));
   MUX2_X1 i_106_0_312 (.A(\mem[71] [7]), .B(data[7]), .S(n_72), .Z(n_106_487));
   MUX2_X1 i_106_0_313 (.A(\mem[71] [6]), .B(data[6]), .S(n_72), .Z(n_106_486));
   MUX2_X1 i_106_0_314 (.A(\mem[71] [5]), .B(data[5]), .S(n_72), .Z(n_106_485));
   MUX2_X1 i_106_0_315 (.A(\mem[71] [4]), .B(data[4]), .S(n_72), .Z(n_106_484));
   MUX2_X1 i_106_0_316 (.A(\mem[71] [3]), .B(data[3]), .S(n_72), .Z(n_106_483));
   MUX2_X1 i_106_0_317 (.A(\mem[71] [2]), .B(data[2]), .S(n_72), .Z(n_106_482));
   MUX2_X1 i_106_0_318 (.A(\mem[71] [1]), .B(data[1]), .S(n_72), .Z(n_106_481));
   MUX2_X1 i_106_0_319 (.A(\mem[71] [0]), .B(data[0]), .S(n_72), .Z(n_106_480));
   MUX2_X1 i_106_0_320 (.A(\mem[72] [15]), .B(data[15]), .S(n_73), .Z(n_106_479));
   MUX2_X1 i_106_0_321 (.A(\mem[72] [14]), .B(data[14]), .S(n_73), .Z(n_106_478));
   MUX2_X1 i_106_0_322 (.A(\mem[72] [13]), .B(data[13]), .S(n_73), .Z(n_106_477));
   MUX2_X1 i_106_0_323 (.A(\mem[72] [12]), .B(data[12]), .S(n_73), .Z(n_106_476));
   MUX2_X1 i_106_0_324 (.A(\mem[72] [11]), .B(data[11]), .S(n_73), .Z(n_106_475));
   MUX2_X1 i_106_0_325 (.A(\mem[72] [10]), .B(data[10]), .S(n_73), .Z(n_106_474));
   MUX2_X1 i_106_0_326 (.A(\mem[72] [9]), .B(data[9]), .S(n_73), .Z(n_106_473));
   MUX2_X1 i_106_0_327 (.A(\mem[72] [8]), .B(data[8]), .S(n_73), .Z(n_106_472));
   MUX2_X1 i_106_0_328 (.A(\mem[72] [7]), .B(data[7]), .S(n_73), .Z(n_106_471));
   MUX2_X1 i_106_0_329 (.A(\mem[72] [6]), .B(data[6]), .S(n_73), .Z(n_106_470));
   MUX2_X1 i_106_0_330 (.A(\mem[72] [5]), .B(data[5]), .S(n_73), .Z(n_106_469));
   MUX2_X1 i_106_0_331 (.A(\mem[72] [4]), .B(data[4]), .S(n_73), .Z(n_106_468));
   MUX2_X1 i_106_0_332 (.A(\mem[72] [3]), .B(data[3]), .S(n_73), .Z(n_106_467));
   MUX2_X1 i_106_0_333 (.A(\mem[72] [2]), .B(data[2]), .S(n_73), .Z(n_106_466));
   MUX2_X1 i_106_0_334 (.A(\mem[72] [1]), .B(data[1]), .S(n_73), .Z(n_106_465));
   MUX2_X1 i_106_0_335 (.A(\mem[72] [0]), .B(data[0]), .S(n_73), .Z(n_106_464));
   MUX2_X1 i_106_0_336 (.A(\mem[73] [15]), .B(data[15]), .S(n_74), .Z(n_106_463));
   MUX2_X1 i_106_0_337 (.A(\mem[73] [14]), .B(data[14]), .S(n_74), .Z(n_106_462));
   MUX2_X1 i_106_0_338 (.A(\mem[73] [13]), .B(data[13]), .S(n_74), .Z(n_106_461));
   MUX2_X1 i_106_0_339 (.A(\mem[73] [12]), .B(data[12]), .S(n_74), .Z(n_106_460));
   MUX2_X1 i_106_0_340 (.A(\mem[73] [11]), .B(data[11]), .S(n_74), .Z(n_106_459));
   MUX2_X1 i_106_0_341 (.A(\mem[73] [10]), .B(data[10]), .S(n_74), .Z(n_106_458));
   MUX2_X1 i_106_0_342 (.A(\mem[73] [9]), .B(data[9]), .S(n_74), .Z(n_106_457));
   MUX2_X1 i_106_0_343 (.A(\mem[73] [8]), .B(data[8]), .S(n_74), .Z(n_106_456));
   MUX2_X1 i_106_0_344 (.A(\mem[73] [7]), .B(data[7]), .S(n_74), .Z(n_106_455));
   MUX2_X1 i_106_0_345 (.A(\mem[73] [6]), .B(data[6]), .S(n_74), .Z(n_106_454));
   MUX2_X1 i_106_0_346 (.A(\mem[73] [5]), .B(data[5]), .S(n_74), .Z(n_106_453));
   MUX2_X1 i_106_0_347 (.A(\mem[73] [4]), .B(data[4]), .S(n_74), .Z(n_106_452));
   MUX2_X1 i_106_0_348 (.A(\mem[73] [3]), .B(data[3]), .S(n_74), .Z(n_106_451));
   MUX2_X1 i_106_0_349 (.A(\mem[73] [2]), .B(data[2]), .S(n_74), .Z(n_106_450));
   MUX2_X1 i_106_0_350 (.A(\mem[73] [1]), .B(data[1]), .S(n_74), .Z(n_106_449));
   MUX2_X1 i_106_0_351 (.A(\mem[73] [0]), .B(data[0]), .S(n_74), .Z(n_106_448));
   MUX2_X1 i_106_0_352 (.A(\mem[74] [15]), .B(data[15]), .S(n_75), .Z(n_106_447));
   MUX2_X1 i_106_0_353 (.A(\mem[74] [14]), .B(data[14]), .S(n_75), .Z(n_106_446));
   MUX2_X1 i_106_0_354 (.A(\mem[74] [13]), .B(data[13]), .S(n_75), .Z(n_106_445));
   MUX2_X1 i_106_0_355 (.A(\mem[74] [12]), .B(data[12]), .S(n_75), .Z(n_106_444));
   MUX2_X1 i_106_0_356 (.A(\mem[74] [11]), .B(data[11]), .S(n_75), .Z(n_106_443));
   MUX2_X1 i_106_0_357 (.A(\mem[74] [10]), .B(data[10]), .S(n_75), .Z(n_106_442));
   MUX2_X1 i_106_0_358 (.A(\mem[74] [9]), .B(data[9]), .S(n_75), .Z(n_106_441));
   MUX2_X1 i_106_0_359 (.A(\mem[74] [8]), .B(data[8]), .S(n_75), .Z(n_106_440));
   MUX2_X1 i_106_0_360 (.A(\mem[74] [7]), .B(data[7]), .S(n_75), .Z(n_106_439));
   MUX2_X1 i_106_0_361 (.A(\mem[74] [6]), .B(data[6]), .S(n_75), .Z(n_106_438));
   MUX2_X1 i_106_0_362 (.A(\mem[74] [5]), .B(data[5]), .S(n_75), .Z(n_106_437));
   MUX2_X1 i_106_0_363 (.A(\mem[74] [4]), .B(data[4]), .S(n_75), .Z(n_106_436));
   MUX2_X1 i_106_0_364 (.A(\mem[74] [3]), .B(data[3]), .S(n_75), .Z(n_106_435));
   MUX2_X1 i_106_0_365 (.A(\mem[74] [2]), .B(data[2]), .S(n_75), .Z(n_106_434));
   MUX2_X1 i_106_0_366 (.A(\mem[74] [1]), .B(data[1]), .S(n_75), .Z(n_106_433));
   MUX2_X1 i_106_0_367 (.A(\mem[74] [0]), .B(data[0]), .S(n_75), .Z(n_106_432));
   MUX2_X1 i_106_0_368 (.A(\mem[75] [15]), .B(data[15]), .S(n_76), .Z(n_106_431));
   MUX2_X1 i_106_0_369 (.A(\mem[75] [14]), .B(data[14]), .S(n_76), .Z(n_106_430));
   MUX2_X1 i_106_0_370 (.A(\mem[75] [13]), .B(data[13]), .S(n_76), .Z(n_106_429));
   MUX2_X1 i_106_0_371 (.A(\mem[75] [12]), .B(data[12]), .S(n_76), .Z(n_106_428));
   MUX2_X1 i_106_0_372 (.A(\mem[75] [11]), .B(data[11]), .S(n_76), .Z(n_106_427));
   MUX2_X1 i_106_0_373 (.A(\mem[75] [10]), .B(data[10]), .S(n_76), .Z(n_106_426));
   MUX2_X1 i_106_0_374 (.A(\mem[75] [9]), .B(data[9]), .S(n_76), .Z(n_106_425));
   MUX2_X1 i_106_0_375 (.A(\mem[75] [8]), .B(data[8]), .S(n_76), .Z(n_106_424));
   MUX2_X1 i_106_0_376 (.A(\mem[75] [7]), .B(data[7]), .S(n_76), .Z(n_106_423));
   MUX2_X1 i_106_0_377 (.A(\mem[75] [6]), .B(data[6]), .S(n_76), .Z(n_106_422));
   MUX2_X1 i_106_0_378 (.A(\mem[75] [5]), .B(data[5]), .S(n_76), .Z(n_106_421));
   MUX2_X1 i_106_0_379 (.A(\mem[75] [4]), .B(data[4]), .S(n_76), .Z(n_106_420));
   MUX2_X1 i_106_0_380 (.A(\mem[75] [3]), .B(data[3]), .S(n_76), .Z(n_106_419));
   MUX2_X1 i_106_0_381 (.A(\mem[75] [2]), .B(data[2]), .S(n_76), .Z(n_106_418));
   MUX2_X1 i_106_0_382 (.A(\mem[75] [1]), .B(data[1]), .S(n_76), .Z(n_106_417));
   MUX2_X1 i_106_0_383 (.A(\mem[75] [0]), .B(data[0]), .S(n_76), .Z(n_106_416));
   MUX2_X1 i_106_0_384 (.A(\mem[76] [15]), .B(data[15]), .S(n_77), .Z(n_106_415));
   MUX2_X1 i_106_0_385 (.A(\mem[76] [14]), .B(data[14]), .S(n_77), .Z(n_106_414));
   MUX2_X1 i_106_0_386 (.A(\mem[76] [13]), .B(data[13]), .S(n_77), .Z(n_106_413));
   MUX2_X1 i_106_0_387 (.A(\mem[76] [12]), .B(data[12]), .S(n_77), .Z(n_106_412));
   MUX2_X1 i_106_0_388 (.A(\mem[76] [11]), .B(data[11]), .S(n_77), .Z(n_106_411));
   MUX2_X1 i_106_0_389 (.A(\mem[76] [10]), .B(data[10]), .S(n_77), .Z(n_106_410));
   MUX2_X1 i_106_0_390 (.A(\mem[76] [9]), .B(data[9]), .S(n_77), .Z(n_106_409));
   MUX2_X1 i_106_0_391 (.A(\mem[76] [8]), .B(data[8]), .S(n_77), .Z(n_106_408));
   MUX2_X1 i_106_0_392 (.A(\mem[76] [7]), .B(data[7]), .S(n_77), .Z(n_106_407));
   MUX2_X1 i_106_0_393 (.A(\mem[76] [6]), .B(data[6]), .S(n_77), .Z(n_106_406));
   MUX2_X1 i_106_0_394 (.A(\mem[76] [5]), .B(data[5]), .S(n_77), .Z(n_106_405));
   MUX2_X1 i_106_0_395 (.A(\mem[76] [4]), .B(data[4]), .S(n_77), .Z(n_106_404));
   MUX2_X1 i_106_0_396 (.A(\mem[76] [3]), .B(data[3]), .S(n_77), .Z(n_106_403));
   MUX2_X1 i_106_0_397 (.A(\mem[76] [2]), .B(data[2]), .S(n_77), .Z(n_106_402));
   MUX2_X1 i_106_0_398 (.A(\mem[76] [1]), .B(data[1]), .S(n_77), .Z(n_106_401));
   MUX2_X1 i_106_0_399 (.A(\mem[76] [0]), .B(data[0]), .S(n_77), .Z(n_106_400));
   MUX2_X1 i_106_0_400 (.A(\mem[77] [15]), .B(data[15]), .S(n_78), .Z(n_106_399));
   MUX2_X1 i_106_0_401 (.A(\mem[77] [14]), .B(data[14]), .S(n_78), .Z(n_106_398));
   MUX2_X1 i_106_0_402 (.A(\mem[77] [13]), .B(data[13]), .S(n_78), .Z(n_106_397));
   MUX2_X1 i_106_0_403 (.A(\mem[77] [12]), .B(data[12]), .S(n_78), .Z(n_106_396));
   MUX2_X1 i_106_0_404 (.A(\mem[77] [11]), .B(data[11]), .S(n_78), .Z(n_106_395));
   MUX2_X1 i_106_0_405 (.A(\mem[77] [10]), .B(data[10]), .S(n_78), .Z(n_106_394));
   MUX2_X1 i_106_0_406 (.A(\mem[77] [9]), .B(data[9]), .S(n_78), .Z(n_106_393));
   MUX2_X1 i_106_0_407 (.A(\mem[77] [8]), .B(data[8]), .S(n_78), .Z(n_106_392));
   MUX2_X1 i_106_0_408 (.A(\mem[77] [7]), .B(data[7]), .S(n_78), .Z(n_106_391));
   MUX2_X1 i_106_0_409 (.A(\mem[77] [6]), .B(data[6]), .S(n_78), .Z(n_106_390));
   MUX2_X1 i_106_0_410 (.A(\mem[77] [5]), .B(data[5]), .S(n_78), .Z(n_106_389));
   MUX2_X1 i_106_0_411 (.A(\mem[77] [4]), .B(data[4]), .S(n_78), .Z(n_106_388));
   MUX2_X1 i_106_0_412 (.A(\mem[77] [3]), .B(data[3]), .S(n_78), .Z(n_106_387));
   MUX2_X1 i_106_0_413 (.A(\mem[77] [2]), .B(data[2]), .S(n_78), .Z(n_106_386));
   MUX2_X1 i_106_0_414 (.A(\mem[77] [1]), .B(data[1]), .S(n_78), .Z(n_106_385));
   MUX2_X1 i_106_0_415 (.A(\mem[77] [0]), .B(data[0]), .S(n_78), .Z(n_106_384));
   MUX2_X1 i_106_0_416 (.A(\mem[78] [15]), .B(data[15]), .S(n_79), .Z(n_106_383));
   MUX2_X1 i_106_0_417 (.A(\mem[78] [14]), .B(data[14]), .S(n_79), .Z(n_106_382));
   MUX2_X1 i_106_0_418 (.A(\mem[78] [13]), .B(data[13]), .S(n_79), .Z(n_106_381));
   MUX2_X1 i_106_0_419 (.A(\mem[78] [12]), .B(data[12]), .S(n_79), .Z(n_106_380));
   MUX2_X1 i_106_0_420 (.A(\mem[78] [11]), .B(data[11]), .S(n_79), .Z(n_106_379));
   MUX2_X1 i_106_0_421 (.A(\mem[78] [10]), .B(data[10]), .S(n_79), .Z(n_106_378));
   MUX2_X1 i_106_0_422 (.A(\mem[78] [9]), .B(data[9]), .S(n_79), .Z(n_106_377));
   MUX2_X1 i_106_0_423 (.A(\mem[78] [8]), .B(data[8]), .S(n_79), .Z(n_106_376));
   MUX2_X1 i_106_0_424 (.A(\mem[78] [7]), .B(data[7]), .S(n_79), .Z(n_106_375));
   MUX2_X1 i_106_0_425 (.A(\mem[78] [6]), .B(data[6]), .S(n_79), .Z(n_106_374));
   MUX2_X1 i_106_0_426 (.A(\mem[78] [5]), .B(data[5]), .S(n_79), .Z(n_106_373));
   MUX2_X1 i_106_0_427 (.A(\mem[78] [4]), .B(data[4]), .S(n_79), .Z(n_106_372));
   MUX2_X1 i_106_0_428 (.A(\mem[78] [3]), .B(data[3]), .S(n_79), .Z(n_106_371));
   MUX2_X1 i_106_0_429 (.A(\mem[78] [2]), .B(data[2]), .S(n_79), .Z(n_106_370));
   MUX2_X1 i_106_0_430 (.A(\mem[78] [1]), .B(data[1]), .S(n_79), .Z(n_106_369));
   MUX2_X1 i_106_0_431 (.A(\mem[78] [0]), .B(data[0]), .S(n_79), .Z(n_106_368));
   MUX2_X1 i_106_0_432 (.A(\mem[79] [15]), .B(data[15]), .S(n_80), .Z(n_106_367));
   MUX2_X1 i_106_0_433 (.A(\mem[79] [14]), .B(data[14]), .S(n_80), .Z(n_106_366));
   MUX2_X1 i_106_0_434 (.A(\mem[79] [13]), .B(data[13]), .S(n_80), .Z(n_106_365));
   MUX2_X1 i_106_0_435 (.A(\mem[79] [12]), .B(data[12]), .S(n_80), .Z(n_106_364));
   MUX2_X1 i_106_0_436 (.A(\mem[79] [11]), .B(data[11]), .S(n_80), .Z(n_106_363));
   MUX2_X1 i_106_0_437 (.A(\mem[79] [10]), .B(data[10]), .S(n_80), .Z(n_106_362));
   MUX2_X1 i_106_0_438 (.A(\mem[79] [9]), .B(data[9]), .S(n_80), .Z(n_106_361));
   MUX2_X1 i_106_0_439 (.A(\mem[79] [8]), .B(data[8]), .S(n_80), .Z(n_106_360));
   MUX2_X1 i_106_0_440 (.A(\mem[79] [7]), .B(data[7]), .S(n_80), .Z(n_106_359));
   MUX2_X1 i_106_0_441 (.A(\mem[79] [6]), .B(data[6]), .S(n_80), .Z(n_106_358));
   MUX2_X1 i_106_0_442 (.A(\mem[79] [5]), .B(data[5]), .S(n_80), .Z(n_106_357));
   MUX2_X1 i_106_0_443 (.A(\mem[79] [4]), .B(data[4]), .S(n_80), .Z(n_106_356));
   MUX2_X1 i_106_0_444 (.A(\mem[79] [3]), .B(data[3]), .S(n_80), .Z(n_106_355));
   MUX2_X1 i_106_0_445 (.A(\mem[79] [2]), .B(data[2]), .S(n_80), .Z(n_106_354));
   MUX2_X1 i_106_0_446 (.A(\mem[79] [1]), .B(data[1]), .S(n_80), .Z(n_106_353));
   MUX2_X1 i_106_0_447 (.A(\mem[79] [0]), .B(data[0]), .S(n_80), .Z(n_106_352));
   MUX2_X1 i_106_0_448 (.A(\mem[80] [15]), .B(data[15]), .S(n_81), .Z(n_106_351));
   MUX2_X1 i_106_0_449 (.A(\mem[80] [14]), .B(data[14]), .S(n_81), .Z(n_106_350));
   MUX2_X1 i_106_0_450 (.A(\mem[80] [13]), .B(data[13]), .S(n_81), .Z(n_106_349));
   MUX2_X1 i_106_0_451 (.A(\mem[80] [12]), .B(data[12]), .S(n_81), .Z(n_106_348));
   MUX2_X1 i_106_0_452 (.A(\mem[80] [11]), .B(data[11]), .S(n_81), .Z(n_106_347));
   MUX2_X1 i_106_0_453 (.A(\mem[80] [10]), .B(data[10]), .S(n_81), .Z(n_106_346));
   MUX2_X1 i_106_0_454 (.A(\mem[80] [9]), .B(data[9]), .S(n_81), .Z(n_106_345));
   MUX2_X1 i_106_0_455 (.A(\mem[80] [8]), .B(data[8]), .S(n_81), .Z(n_106_344));
   MUX2_X1 i_106_0_456 (.A(\mem[80] [7]), .B(data[7]), .S(n_81), .Z(n_106_343));
   MUX2_X1 i_106_0_457 (.A(\mem[80] [6]), .B(data[6]), .S(n_81), .Z(n_106_342));
   MUX2_X1 i_106_0_458 (.A(\mem[80] [5]), .B(data[5]), .S(n_81), .Z(n_106_341));
   MUX2_X1 i_106_0_459 (.A(\mem[80] [4]), .B(data[4]), .S(n_81), .Z(n_106_340));
   MUX2_X1 i_106_0_460 (.A(\mem[80] [3]), .B(data[3]), .S(n_81), .Z(n_106_339));
   MUX2_X1 i_106_0_461 (.A(\mem[80] [2]), .B(data[2]), .S(n_81), .Z(n_106_338));
   MUX2_X1 i_106_0_462 (.A(\mem[80] [1]), .B(data[1]), .S(n_81), .Z(n_106_337));
   MUX2_X1 i_106_0_463 (.A(\mem[80] [0]), .B(data[0]), .S(n_81), .Z(n_106_336));
   MUX2_X1 i_106_0_464 (.A(\mem[81] [15]), .B(data[15]), .S(n_82), .Z(n_106_335));
   MUX2_X1 i_106_0_465 (.A(\mem[81] [14]), .B(data[14]), .S(n_82), .Z(n_106_334));
   MUX2_X1 i_106_0_466 (.A(\mem[81] [13]), .B(data[13]), .S(n_82), .Z(n_106_333));
   MUX2_X1 i_106_0_467 (.A(\mem[81] [12]), .B(data[12]), .S(n_82), .Z(n_106_332));
   MUX2_X1 i_106_0_468 (.A(\mem[81] [11]), .B(data[11]), .S(n_82), .Z(n_106_331));
   MUX2_X1 i_106_0_469 (.A(\mem[81] [10]), .B(data[10]), .S(n_82), .Z(n_106_330));
   MUX2_X1 i_106_0_470 (.A(\mem[81] [9]), .B(data[9]), .S(n_82), .Z(n_106_329));
   MUX2_X1 i_106_0_471 (.A(\mem[81] [8]), .B(data[8]), .S(n_82), .Z(n_106_328));
   MUX2_X1 i_106_0_472 (.A(\mem[81] [7]), .B(data[7]), .S(n_82), .Z(n_106_327));
   MUX2_X1 i_106_0_473 (.A(\mem[81] [6]), .B(data[6]), .S(n_82), .Z(n_106_326));
   MUX2_X1 i_106_0_474 (.A(\mem[81] [5]), .B(data[5]), .S(n_82), .Z(n_106_325));
   MUX2_X1 i_106_0_475 (.A(\mem[81] [4]), .B(data[4]), .S(n_82), .Z(n_106_324));
   MUX2_X1 i_106_0_476 (.A(\mem[81] [3]), .B(data[3]), .S(n_82), .Z(n_106_323));
   MUX2_X1 i_106_0_477 (.A(\mem[81] [2]), .B(data[2]), .S(n_82), .Z(n_106_322));
   MUX2_X1 i_106_0_478 (.A(\mem[81] [1]), .B(data[1]), .S(n_82), .Z(n_106_321));
   MUX2_X1 i_106_0_479 (.A(\mem[81] [0]), .B(data[0]), .S(n_82), .Z(n_106_320));
   MUX2_X1 i_106_0_480 (.A(\mem[82] [15]), .B(data[15]), .S(n_83), .Z(n_106_319));
   MUX2_X1 i_106_0_481 (.A(\mem[82] [14]), .B(data[14]), .S(n_83), .Z(n_106_318));
   MUX2_X1 i_106_0_482 (.A(\mem[82] [13]), .B(data[13]), .S(n_83), .Z(n_106_317));
   MUX2_X1 i_106_0_483 (.A(\mem[82] [12]), .B(data[12]), .S(n_83), .Z(n_106_316));
   MUX2_X1 i_106_0_484 (.A(\mem[82] [11]), .B(data[11]), .S(n_83), .Z(n_106_315));
   MUX2_X1 i_106_0_485 (.A(\mem[82] [10]), .B(data[10]), .S(n_83), .Z(n_106_314));
   MUX2_X1 i_106_0_486 (.A(\mem[82] [9]), .B(data[9]), .S(n_83), .Z(n_106_313));
   MUX2_X1 i_106_0_487 (.A(\mem[82] [8]), .B(data[8]), .S(n_83), .Z(n_106_312));
   MUX2_X1 i_106_0_488 (.A(\mem[82] [7]), .B(data[7]), .S(n_83), .Z(n_106_311));
   MUX2_X1 i_106_0_489 (.A(\mem[82] [6]), .B(data[6]), .S(n_83), .Z(n_106_310));
   MUX2_X1 i_106_0_490 (.A(\mem[82] [5]), .B(data[5]), .S(n_83), .Z(n_106_309));
   MUX2_X1 i_106_0_491 (.A(\mem[82] [4]), .B(data[4]), .S(n_83), .Z(n_106_308));
   MUX2_X1 i_106_0_492 (.A(\mem[82] [3]), .B(data[3]), .S(n_83), .Z(n_106_307));
   MUX2_X1 i_106_0_493 (.A(\mem[82] [2]), .B(data[2]), .S(n_83), .Z(n_106_306));
   MUX2_X1 i_106_0_494 (.A(\mem[82] [1]), .B(data[1]), .S(n_83), .Z(n_106_305));
   MUX2_X1 i_106_0_495 (.A(\mem[82] [0]), .B(data[0]), .S(n_83), .Z(n_106_304));
   MUX2_X1 i_106_0_496 (.A(\mem[83] [15]), .B(data[15]), .S(n_84), .Z(n_106_303));
   MUX2_X1 i_106_0_497 (.A(\mem[83] [14]), .B(data[14]), .S(n_84), .Z(n_106_302));
   MUX2_X1 i_106_0_498 (.A(\mem[83] [13]), .B(data[13]), .S(n_84), .Z(n_106_301));
   MUX2_X1 i_106_0_499 (.A(\mem[83] [12]), .B(data[12]), .S(n_84), .Z(n_106_300));
   MUX2_X1 i_106_0_500 (.A(\mem[83] [11]), .B(data[11]), .S(n_84), .Z(n_106_299));
   MUX2_X1 i_106_0_501 (.A(\mem[83] [10]), .B(data[10]), .S(n_84), .Z(n_106_298));
   MUX2_X1 i_106_0_502 (.A(\mem[83] [9]), .B(data[9]), .S(n_84), .Z(n_106_297));
   MUX2_X1 i_106_0_503 (.A(\mem[83] [8]), .B(data[8]), .S(n_84), .Z(n_106_296));
   MUX2_X1 i_106_0_504 (.A(\mem[83] [7]), .B(data[7]), .S(n_84), .Z(n_106_295));
   MUX2_X1 i_106_0_505 (.A(\mem[83] [6]), .B(data[6]), .S(n_84), .Z(n_106_294));
   MUX2_X1 i_106_0_506 (.A(\mem[83] [5]), .B(data[5]), .S(n_84), .Z(n_106_293));
   MUX2_X1 i_106_0_507 (.A(\mem[83] [4]), .B(data[4]), .S(n_84), .Z(n_106_292));
   MUX2_X1 i_106_0_508 (.A(\mem[83] [3]), .B(data[3]), .S(n_84), .Z(n_106_291));
   MUX2_X1 i_106_0_509 (.A(\mem[83] [2]), .B(data[2]), .S(n_84), .Z(n_106_290));
   MUX2_X1 i_106_0_510 (.A(\mem[83] [1]), .B(data[1]), .S(n_84), .Z(n_106_289));
   MUX2_X1 i_106_0_511 (.A(\mem[83] [0]), .B(data[0]), .S(n_84), .Z(n_106_288));
   MUX2_X1 i_106_0_512 (.A(\mem[84] [15]), .B(data[15]), .S(n_85), .Z(n_106_287));
   MUX2_X1 i_106_0_513 (.A(\mem[84] [14]), .B(data[14]), .S(n_85), .Z(n_106_286));
   MUX2_X1 i_106_0_514 (.A(\mem[84] [13]), .B(data[13]), .S(n_85), .Z(n_106_285));
   MUX2_X1 i_106_0_515 (.A(\mem[84] [12]), .B(data[12]), .S(n_85), .Z(n_106_284));
   MUX2_X1 i_106_0_516 (.A(\mem[84] [11]), .B(data[11]), .S(n_85), .Z(n_106_283));
   MUX2_X1 i_106_0_517 (.A(\mem[84] [10]), .B(data[10]), .S(n_85), .Z(n_106_282));
   MUX2_X1 i_106_0_518 (.A(\mem[84] [9]), .B(data[9]), .S(n_85), .Z(n_106_281));
   MUX2_X1 i_106_0_519 (.A(\mem[84] [8]), .B(data[8]), .S(n_85), .Z(n_106_280));
   MUX2_X1 i_106_0_520 (.A(\mem[84] [7]), .B(data[7]), .S(n_85), .Z(n_106_279));
   MUX2_X1 i_106_0_521 (.A(\mem[84] [6]), .B(data[6]), .S(n_85), .Z(n_106_278));
   MUX2_X1 i_106_0_522 (.A(\mem[84] [5]), .B(data[5]), .S(n_85), .Z(n_106_277));
   MUX2_X1 i_106_0_523 (.A(\mem[84] [4]), .B(data[4]), .S(n_85), .Z(n_106_276));
   MUX2_X1 i_106_0_524 (.A(\mem[84] [3]), .B(data[3]), .S(n_85), .Z(n_106_275));
   MUX2_X1 i_106_0_525 (.A(\mem[84] [2]), .B(data[2]), .S(n_85), .Z(n_106_274));
   MUX2_X1 i_106_0_526 (.A(\mem[84] [1]), .B(data[1]), .S(n_85), .Z(n_106_273));
   MUX2_X1 i_106_0_527 (.A(\mem[84] [0]), .B(data[0]), .S(n_85), .Z(n_106_272));
   MUX2_X1 i_106_0_528 (.A(\mem[85] [15]), .B(data[15]), .S(n_86), .Z(n_106_271));
   MUX2_X1 i_106_0_529 (.A(\mem[85] [14]), .B(data[14]), .S(n_86), .Z(n_106_270));
   MUX2_X1 i_106_0_530 (.A(\mem[85] [13]), .B(data[13]), .S(n_86), .Z(n_106_269));
   MUX2_X1 i_106_0_531 (.A(\mem[85] [12]), .B(data[12]), .S(n_86), .Z(n_106_268));
   MUX2_X1 i_106_0_532 (.A(\mem[85] [11]), .B(data[11]), .S(n_86), .Z(n_106_267));
   MUX2_X1 i_106_0_533 (.A(\mem[85] [10]), .B(data[10]), .S(n_86), .Z(n_106_266));
   MUX2_X1 i_106_0_534 (.A(\mem[85] [9]), .B(data[9]), .S(n_86), .Z(n_106_265));
   MUX2_X1 i_106_0_535 (.A(\mem[85] [8]), .B(data[8]), .S(n_86), .Z(n_106_264));
   MUX2_X1 i_106_0_536 (.A(\mem[85] [7]), .B(data[7]), .S(n_86), .Z(n_106_263));
   MUX2_X1 i_106_0_537 (.A(\mem[85] [6]), .B(data[6]), .S(n_86), .Z(n_106_262));
   MUX2_X1 i_106_0_538 (.A(\mem[85] [5]), .B(data[5]), .S(n_86), .Z(n_106_261));
   MUX2_X1 i_106_0_539 (.A(\mem[85] [4]), .B(data[4]), .S(n_86), .Z(n_106_260));
   MUX2_X1 i_106_0_540 (.A(\mem[85] [3]), .B(data[3]), .S(n_86), .Z(n_106_259));
   MUX2_X1 i_106_0_541 (.A(\mem[85] [2]), .B(data[2]), .S(n_86), .Z(n_106_258));
   MUX2_X1 i_106_0_542 (.A(\mem[85] [1]), .B(data[1]), .S(n_86), .Z(n_106_257));
   MUX2_X1 i_106_0_543 (.A(\mem[85] [0]), .B(data[0]), .S(n_86), .Z(n_106_256));
   MUX2_X1 i_106_0_544 (.A(\mem[86] [15]), .B(data[15]), .S(n_87), .Z(n_106_255));
   MUX2_X1 i_106_0_545 (.A(\mem[86] [14]), .B(data[14]), .S(n_87), .Z(n_106_254));
   MUX2_X1 i_106_0_546 (.A(\mem[86] [13]), .B(data[13]), .S(n_87), .Z(n_106_253));
   MUX2_X1 i_106_0_547 (.A(\mem[86] [12]), .B(data[12]), .S(n_87), .Z(n_106_252));
   MUX2_X1 i_106_0_548 (.A(\mem[86] [11]), .B(data[11]), .S(n_87), .Z(n_106_251));
   MUX2_X1 i_106_0_549 (.A(\mem[86] [10]), .B(data[10]), .S(n_87), .Z(n_106_250));
   MUX2_X1 i_106_0_550 (.A(\mem[86] [9]), .B(data[9]), .S(n_87), .Z(n_106_249));
   MUX2_X1 i_106_0_551 (.A(\mem[86] [8]), .B(data[8]), .S(n_87), .Z(n_106_248));
   MUX2_X1 i_106_0_552 (.A(\mem[86] [7]), .B(data[7]), .S(n_87), .Z(n_106_247));
   MUX2_X1 i_106_0_553 (.A(\mem[86] [6]), .B(data[6]), .S(n_87), .Z(n_106_246));
   MUX2_X1 i_106_0_554 (.A(\mem[86] [5]), .B(data[5]), .S(n_87), .Z(n_106_245));
   MUX2_X1 i_106_0_555 (.A(\mem[86] [4]), .B(data[4]), .S(n_87), .Z(n_106_244));
   MUX2_X1 i_106_0_556 (.A(\mem[86] [3]), .B(data[3]), .S(n_87), .Z(n_106_243));
   MUX2_X1 i_106_0_557 (.A(\mem[86] [2]), .B(data[2]), .S(n_87), .Z(n_106_242));
   MUX2_X1 i_106_0_558 (.A(\mem[86] [1]), .B(data[1]), .S(n_87), .Z(n_106_241));
   MUX2_X1 i_106_0_559 (.A(\mem[86] [0]), .B(data[0]), .S(n_87), .Z(n_106_240));
   MUX2_X1 i_106_0_560 (.A(\mem[87] [15]), .B(data[15]), .S(n_88), .Z(n_106_239));
   MUX2_X1 i_106_0_561 (.A(\mem[87] [14]), .B(data[14]), .S(n_88), .Z(n_106_238));
   MUX2_X1 i_106_0_562 (.A(\mem[87] [13]), .B(data[13]), .S(n_88), .Z(n_106_237));
   MUX2_X1 i_106_0_563 (.A(\mem[87] [12]), .B(data[12]), .S(n_88), .Z(n_106_236));
   MUX2_X1 i_106_0_564 (.A(\mem[87] [11]), .B(data[11]), .S(n_88), .Z(n_106_235));
   MUX2_X1 i_106_0_565 (.A(\mem[87] [10]), .B(data[10]), .S(n_88), .Z(n_106_234));
   MUX2_X1 i_106_0_566 (.A(\mem[87] [9]), .B(data[9]), .S(n_88), .Z(n_106_233));
   MUX2_X1 i_106_0_567 (.A(\mem[87] [8]), .B(data[8]), .S(n_88), .Z(n_106_232));
   MUX2_X1 i_106_0_568 (.A(\mem[87] [7]), .B(data[7]), .S(n_88), .Z(n_106_231));
   MUX2_X1 i_106_0_569 (.A(\mem[87] [6]), .B(data[6]), .S(n_88), .Z(n_106_230));
   MUX2_X1 i_106_0_570 (.A(\mem[87] [5]), .B(data[5]), .S(n_88), .Z(n_106_229));
   MUX2_X1 i_106_0_571 (.A(\mem[87] [4]), .B(data[4]), .S(n_88), .Z(n_106_228));
   MUX2_X1 i_106_0_572 (.A(\mem[87] [3]), .B(data[3]), .S(n_88), .Z(n_106_227));
   MUX2_X1 i_106_0_573 (.A(\mem[87] [2]), .B(data[2]), .S(n_88), .Z(n_106_226));
   MUX2_X1 i_106_0_574 (.A(\mem[87] [1]), .B(data[1]), .S(n_88), .Z(n_106_225));
   MUX2_X1 i_106_0_575 (.A(\mem[87] [0]), .B(data[0]), .S(n_88), .Z(n_106_224));
   MUX2_X1 i_106_0_576 (.A(\mem[88] [15]), .B(data[15]), .S(n_89), .Z(n_106_223));
   MUX2_X1 i_106_0_577 (.A(\mem[88] [14]), .B(data[14]), .S(n_89), .Z(n_106_222));
   MUX2_X1 i_106_0_578 (.A(\mem[88] [13]), .B(data[13]), .S(n_89), .Z(n_106_221));
   MUX2_X1 i_106_0_579 (.A(\mem[88] [12]), .B(data[12]), .S(n_89), .Z(n_106_220));
   MUX2_X1 i_106_0_580 (.A(\mem[88] [11]), .B(data[11]), .S(n_89), .Z(n_106_219));
   MUX2_X1 i_106_0_581 (.A(\mem[88] [10]), .B(data[10]), .S(n_89), .Z(n_106_218));
   MUX2_X1 i_106_0_582 (.A(\mem[88] [9]), .B(data[9]), .S(n_89), .Z(n_106_217));
   MUX2_X1 i_106_0_583 (.A(\mem[88] [8]), .B(data[8]), .S(n_89), .Z(n_106_216));
   MUX2_X1 i_106_0_584 (.A(\mem[88] [7]), .B(data[7]), .S(n_89), .Z(n_106_215));
   MUX2_X1 i_106_0_585 (.A(\mem[88] [6]), .B(data[6]), .S(n_89), .Z(n_106_214));
   MUX2_X1 i_106_0_586 (.A(\mem[88] [5]), .B(data[5]), .S(n_89), .Z(n_106_213));
   MUX2_X1 i_106_0_587 (.A(\mem[88] [4]), .B(data[4]), .S(n_89), .Z(n_106_212));
   MUX2_X1 i_106_0_588 (.A(\mem[88] [3]), .B(data[3]), .S(n_89), .Z(n_106_211));
   MUX2_X1 i_106_0_589 (.A(\mem[88] [2]), .B(data[2]), .S(n_89), .Z(n_106_210));
   MUX2_X1 i_106_0_590 (.A(\mem[88] [1]), .B(data[1]), .S(n_89), .Z(n_106_209));
   MUX2_X1 i_106_0_591 (.A(\mem[88] [0]), .B(data[0]), .S(n_89), .Z(n_106_208));
   MUX2_X1 i_106_0_592 (.A(\mem[89] [15]), .B(data[15]), .S(n_90), .Z(n_106_207));
   MUX2_X1 i_106_0_593 (.A(\mem[89] [14]), .B(data[14]), .S(n_90), .Z(n_106_206));
   MUX2_X1 i_106_0_594 (.A(\mem[89] [13]), .B(data[13]), .S(n_90), .Z(n_106_205));
   MUX2_X1 i_106_0_595 (.A(\mem[89] [12]), .B(data[12]), .S(n_90), .Z(n_106_204));
   MUX2_X1 i_106_0_596 (.A(\mem[89] [11]), .B(data[11]), .S(n_90), .Z(n_106_203));
   MUX2_X1 i_106_0_597 (.A(\mem[89] [10]), .B(data[10]), .S(n_90), .Z(n_106_202));
   MUX2_X1 i_106_0_598 (.A(\mem[89] [9]), .B(data[9]), .S(n_90), .Z(n_106_201));
   MUX2_X1 i_106_0_599 (.A(\mem[89] [8]), .B(data[8]), .S(n_90), .Z(n_106_200));
   MUX2_X1 i_106_0_600 (.A(\mem[89] [7]), .B(data[7]), .S(n_90), .Z(n_106_199));
   MUX2_X1 i_106_0_601 (.A(\mem[89] [6]), .B(data[6]), .S(n_90), .Z(n_106_198));
   MUX2_X1 i_106_0_602 (.A(\mem[89] [5]), .B(data[5]), .S(n_90), .Z(n_106_197));
   MUX2_X1 i_106_0_603 (.A(\mem[89] [4]), .B(data[4]), .S(n_90), .Z(n_106_196));
   MUX2_X1 i_106_0_604 (.A(\mem[89] [3]), .B(data[3]), .S(n_90), .Z(n_106_195));
   MUX2_X1 i_106_0_605 (.A(\mem[89] [2]), .B(data[2]), .S(n_90), .Z(n_106_194));
   MUX2_X1 i_106_0_606 (.A(\mem[89] [1]), .B(data[1]), .S(n_90), .Z(n_106_193));
   MUX2_X1 i_106_0_607 (.A(\mem[89] [0]), .B(data[0]), .S(n_90), .Z(n_106_192));
   MUX2_X1 i_106_0_608 (.A(\mem[90] [15]), .B(data[15]), .S(n_91), .Z(n_106_191));
   MUX2_X1 i_106_0_609 (.A(\mem[90] [14]), .B(data[14]), .S(n_91), .Z(n_106_190));
   MUX2_X1 i_106_0_610 (.A(\mem[90] [13]), .B(data[13]), .S(n_91), .Z(n_106_189));
   MUX2_X1 i_106_0_611 (.A(\mem[90] [12]), .B(data[12]), .S(n_91), .Z(n_106_188));
   MUX2_X1 i_106_0_612 (.A(\mem[90] [11]), .B(data[11]), .S(n_91), .Z(n_106_187));
   MUX2_X1 i_106_0_613 (.A(\mem[90] [10]), .B(data[10]), .S(n_91), .Z(n_106_186));
   MUX2_X1 i_106_0_614 (.A(\mem[90] [9]), .B(data[9]), .S(n_91), .Z(n_106_185));
   MUX2_X1 i_106_0_615 (.A(\mem[90] [8]), .B(data[8]), .S(n_91), .Z(n_106_184));
   MUX2_X1 i_106_0_616 (.A(\mem[90] [7]), .B(data[7]), .S(n_91), .Z(n_106_183));
   MUX2_X1 i_106_0_617 (.A(\mem[90] [6]), .B(data[6]), .S(n_91), .Z(n_106_182));
   MUX2_X1 i_106_0_618 (.A(\mem[90] [5]), .B(data[5]), .S(n_91), .Z(n_106_181));
   MUX2_X1 i_106_0_619 (.A(\mem[90] [4]), .B(data[4]), .S(n_91), .Z(n_106_180));
   MUX2_X1 i_106_0_620 (.A(\mem[90] [3]), .B(data[3]), .S(n_91), .Z(n_106_179));
   MUX2_X1 i_106_0_621 (.A(\mem[90] [2]), .B(data[2]), .S(n_91), .Z(n_106_178));
   MUX2_X1 i_106_0_622 (.A(\mem[90] [1]), .B(data[1]), .S(n_91), .Z(n_106_177));
   MUX2_X1 i_106_0_623 (.A(\mem[90] [0]), .B(data[0]), .S(n_91), .Z(n_106_176));
   MUX2_X1 i_106_0_624 (.A(\mem[91] [15]), .B(data[15]), .S(n_92), .Z(n_106_175));
   MUX2_X1 i_106_0_625 (.A(\mem[91] [14]), .B(data[14]), .S(n_92), .Z(n_106_174));
   MUX2_X1 i_106_0_626 (.A(\mem[91] [13]), .B(data[13]), .S(n_92), .Z(n_106_173));
   MUX2_X1 i_106_0_627 (.A(\mem[91] [12]), .B(data[12]), .S(n_92), .Z(n_106_172));
   MUX2_X1 i_106_0_628 (.A(\mem[91] [11]), .B(data[11]), .S(n_92), .Z(n_106_171));
   MUX2_X1 i_106_0_629 (.A(\mem[91] [10]), .B(data[10]), .S(n_92), .Z(n_106_170));
   MUX2_X1 i_106_0_630 (.A(\mem[91] [9]), .B(data[9]), .S(n_92), .Z(n_106_169));
   MUX2_X1 i_106_0_631 (.A(\mem[91] [8]), .B(data[8]), .S(n_92), .Z(n_106_168));
   MUX2_X1 i_106_0_632 (.A(\mem[91] [7]), .B(data[7]), .S(n_92), .Z(n_106_167));
   MUX2_X1 i_106_0_633 (.A(\mem[91] [6]), .B(data[6]), .S(n_92), .Z(n_106_166));
   MUX2_X1 i_106_0_634 (.A(\mem[91] [5]), .B(data[5]), .S(n_92), .Z(n_106_165));
   MUX2_X1 i_106_0_635 (.A(\mem[91] [4]), .B(data[4]), .S(n_92), .Z(n_106_164));
   MUX2_X1 i_106_0_636 (.A(\mem[91] [3]), .B(data[3]), .S(n_92), .Z(n_106_163));
   MUX2_X1 i_106_0_637 (.A(\mem[91] [2]), .B(data[2]), .S(n_92), .Z(n_106_162));
   MUX2_X1 i_106_0_638 (.A(\mem[91] [1]), .B(data[1]), .S(n_92), .Z(n_106_161));
   MUX2_X1 i_106_0_639 (.A(\mem[91] [0]), .B(data[0]), .S(n_92), .Z(n_106_160));
   MUX2_X1 i_106_0_640 (.A(\mem[92] [15]), .B(data[15]), .S(n_93), .Z(n_106_159));
   MUX2_X1 i_106_0_641 (.A(\mem[92] [14]), .B(data[14]), .S(n_93), .Z(n_106_158));
   MUX2_X1 i_106_0_642 (.A(\mem[92] [13]), .B(data[13]), .S(n_93), .Z(n_106_157));
   MUX2_X1 i_106_0_643 (.A(\mem[92] [12]), .B(data[12]), .S(n_93), .Z(n_106_156));
   MUX2_X1 i_106_0_644 (.A(\mem[92] [11]), .B(data[11]), .S(n_93), .Z(n_106_155));
   MUX2_X1 i_106_0_645 (.A(\mem[92] [10]), .B(data[10]), .S(n_93), .Z(n_106_154));
   MUX2_X1 i_106_0_646 (.A(\mem[92] [9]), .B(data[9]), .S(n_93), .Z(n_106_153));
   MUX2_X1 i_106_0_647 (.A(\mem[92] [8]), .B(data[8]), .S(n_93), .Z(n_106_152));
   MUX2_X1 i_106_0_648 (.A(\mem[92] [7]), .B(data[7]), .S(n_93), .Z(n_106_151));
   MUX2_X1 i_106_0_649 (.A(\mem[92] [6]), .B(data[6]), .S(n_93), .Z(n_106_150));
   MUX2_X1 i_106_0_650 (.A(\mem[92] [5]), .B(data[5]), .S(n_93), .Z(n_106_149));
   MUX2_X1 i_106_0_651 (.A(\mem[92] [4]), .B(data[4]), .S(n_93), .Z(n_106_148));
   MUX2_X1 i_106_0_652 (.A(\mem[92] [3]), .B(data[3]), .S(n_93), .Z(n_106_147));
   MUX2_X1 i_106_0_653 (.A(\mem[92] [2]), .B(data[2]), .S(n_93), .Z(n_106_146));
   MUX2_X1 i_106_0_654 (.A(\mem[92] [1]), .B(data[1]), .S(n_93), .Z(n_106_145));
   MUX2_X1 i_106_0_655 (.A(\mem[92] [0]), .B(data[0]), .S(n_93), .Z(n_106_144));
   MUX2_X1 i_106_0_656 (.A(\mem[93] [15]), .B(data[15]), .S(n_94), .Z(n_106_143));
   MUX2_X1 i_106_0_657 (.A(\mem[93] [14]), .B(data[14]), .S(n_94), .Z(n_106_142));
   MUX2_X1 i_106_0_658 (.A(\mem[93] [13]), .B(data[13]), .S(n_94), .Z(n_106_141));
   MUX2_X1 i_106_0_659 (.A(\mem[93] [12]), .B(data[12]), .S(n_94), .Z(n_106_140));
   MUX2_X1 i_106_0_660 (.A(\mem[93] [11]), .B(data[11]), .S(n_94), .Z(n_106_139));
   MUX2_X1 i_106_0_661 (.A(\mem[93] [10]), .B(data[10]), .S(n_94), .Z(n_106_138));
   MUX2_X1 i_106_0_662 (.A(\mem[93] [9]), .B(data[9]), .S(n_94), .Z(n_106_137));
   MUX2_X1 i_106_0_663 (.A(\mem[93] [8]), .B(data[8]), .S(n_94), .Z(n_106_136));
   MUX2_X1 i_106_0_664 (.A(\mem[93] [7]), .B(data[7]), .S(n_94), .Z(n_106_135));
   MUX2_X1 i_106_0_665 (.A(\mem[93] [6]), .B(data[6]), .S(n_94), .Z(n_106_134));
   MUX2_X1 i_106_0_666 (.A(\mem[93] [5]), .B(data[5]), .S(n_94), .Z(n_106_133));
   MUX2_X1 i_106_0_667 (.A(\mem[93] [4]), .B(data[4]), .S(n_94), .Z(n_106_132));
   MUX2_X1 i_106_0_668 (.A(\mem[93] [3]), .B(data[3]), .S(n_94), .Z(n_106_131));
   MUX2_X1 i_106_0_669 (.A(\mem[93] [2]), .B(data[2]), .S(n_94), .Z(n_106_130));
   MUX2_X1 i_106_0_670 (.A(\mem[93] [1]), .B(data[1]), .S(n_94), .Z(n_106_129));
   MUX2_X1 i_106_0_671 (.A(\mem[93] [0]), .B(data[0]), .S(n_94), .Z(n_106_128));
   MUX2_X1 i_106_0_672 (.A(\mem[94] [15]), .B(data[15]), .S(n_95), .Z(n_106_127));
   MUX2_X1 i_106_0_673 (.A(\mem[94] [14]), .B(data[14]), .S(n_95), .Z(n_106_126));
   MUX2_X1 i_106_0_674 (.A(\mem[94] [13]), .B(data[13]), .S(n_95), .Z(n_106_125));
   MUX2_X1 i_106_0_675 (.A(\mem[94] [12]), .B(data[12]), .S(n_95), .Z(n_106_124));
   MUX2_X1 i_106_0_676 (.A(\mem[94] [11]), .B(data[11]), .S(n_95), .Z(n_106_123));
   MUX2_X1 i_106_0_677 (.A(\mem[94] [10]), .B(data[10]), .S(n_95), .Z(n_106_122));
   MUX2_X1 i_106_0_678 (.A(\mem[94] [9]), .B(data[9]), .S(n_95), .Z(n_106_121));
   MUX2_X1 i_106_0_679 (.A(\mem[94] [8]), .B(data[8]), .S(n_95), .Z(n_106_120));
   MUX2_X1 i_106_0_680 (.A(\mem[94] [7]), .B(data[7]), .S(n_95), .Z(n_106_119));
   MUX2_X1 i_106_0_681 (.A(\mem[94] [6]), .B(data[6]), .S(n_95), .Z(n_106_118));
   MUX2_X1 i_106_0_682 (.A(\mem[94] [5]), .B(data[5]), .S(n_95), .Z(n_106_117));
   MUX2_X1 i_106_0_683 (.A(\mem[94] [4]), .B(data[4]), .S(n_95), .Z(n_106_116));
   MUX2_X1 i_106_0_684 (.A(\mem[94] [3]), .B(data[3]), .S(n_95), .Z(n_106_115));
   MUX2_X1 i_106_0_685 (.A(\mem[94] [2]), .B(data[2]), .S(n_95), .Z(n_106_114));
   MUX2_X1 i_106_0_686 (.A(\mem[94] [1]), .B(data[1]), .S(n_95), .Z(n_106_113));
   MUX2_X1 i_106_0_687 (.A(\mem[94] [0]), .B(data[0]), .S(n_95), .Z(n_106_112));
   MUX2_X1 i_106_0_688 (.A(\mem[95] [15]), .B(data[15]), .S(n_96), .Z(n_106_111));
   MUX2_X1 i_106_0_689 (.A(\mem[95] [14]), .B(data[14]), .S(n_96), .Z(n_106_110));
   MUX2_X1 i_106_0_690 (.A(\mem[95] [13]), .B(data[13]), .S(n_96), .Z(n_106_109));
   MUX2_X1 i_106_0_691 (.A(\mem[95] [12]), .B(data[12]), .S(n_96), .Z(n_106_108));
   MUX2_X1 i_106_0_692 (.A(\mem[95] [11]), .B(data[11]), .S(n_96), .Z(n_106_107));
   MUX2_X1 i_106_0_693 (.A(\mem[95] [10]), .B(data[10]), .S(n_96), .Z(n_106_106));
   MUX2_X1 i_106_0_694 (.A(\mem[95] [9]), .B(data[9]), .S(n_96), .Z(n_106_105));
   MUX2_X1 i_106_0_695 (.A(\mem[95] [8]), .B(data[8]), .S(n_96), .Z(n_106_104));
   MUX2_X1 i_106_0_696 (.A(\mem[95] [7]), .B(data[7]), .S(n_96), .Z(n_106_103));
   MUX2_X1 i_106_0_697 (.A(\mem[95] [6]), .B(data[6]), .S(n_96), .Z(n_106_102));
   MUX2_X1 i_106_0_698 (.A(\mem[95] [5]), .B(data[5]), .S(n_96), .Z(n_106_101));
   MUX2_X1 i_106_0_699 (.A(\mem[95] [4]), .B(data[4]), .S(n_96), .Z(n_106_100));
   MUX2_X1 i_106_0_700 (.A(\mem[95] [3]), .B(data[3]), .S(n_96), .Z(n_106_99));
   MUX2_X1 i_106_0_701 (.A(\mem[95] [2]), .B(data[2]), .S(n_96), .Z(n_106_98));
   MUX2_X1 i_106_0_702 (.A(\mem[95] [1]), .B(data[1]), .S(n_96), .Z(n_106_97));
   MUX2_X1 i_106_0_703 (.A(\mem[95] [0]), .B(data[0]), .S(n_96), .Z(n_106_96));
   MUX2_X1 i_106_0_704 (.A(\mem[96] [15]), .B(data[15]), .S(n_97), .Z(n_106_95));
   MUX2_X1 i_106_0_705 (.A(\mem[96] [14]), .B(data[14]), .S(n_97), .Z(n_106_94));
   MUX2_X1 i_106_0_706 (.A(\mem[96] [13]), .B(data[13]), .S(n_97), .Z(n_106_93));
   MUX2_X1 i_106_0_707 (.A(\mem[96] [12]), .B(data[12]), .S(n_97), .Z(n_106_92));
   MUX2_X1 i_106_0_708 (.A(\mem[96] [11]), .B(data[11]), .S(n_97), .Z(n_106_91));
   MUX2_X1 i_106_0_709 (.A(\mem[96] [10]), .B(data[10]), .S(n_97), .Z(n_106_90));
   MUX2_X1 i_106_0_710 (.A(\mem[96] [9]), .B(data[9]), .S(n_97), .Z(n_106_89));
   MUX2_X1 i_106_0_711 (.A(\mem[96] [8]), .B(data[8]), .S(n_97), .Z(n_106_88));
   MUX2_X1 i_106_0_712 (.A(\mem[96] [7]), .B(data[7]), .S(n_97), .Z(n_106_87));
   MUX2_X1 i_106_0_713 (.A(\mem[96] [6]), .B(data[6]), .S(n_97), .Z(n_106_86));
   MUX2_X1 i_106_0_714 (.A(\mem[96] [5]), .B(data[5]), .S(n_97), .Z(n_106_85));
   MUX2_X1 i_106_0_715 (.A(\mem[96] [4]), .B(data[4]), .S(n_97), .Z(n_106_84));
   MUX2_X1 i_106_0_716 (.A(\mem[96] [3]), .B(data[3]), .S(n_97), .Z(n_106_83));
   MUX2_X1 i_106_0_717 (.A(\mem[96] [2]), .B(data[2]), .S(n_97), .Z(n_106_82));
   MUX2_X1 i_106_0_718 (.A(\mem[96] [1]), .B(data[1]), .S(n_97), .Z(n_106_81));
   MUX2_X1 i_106_0_719 (.A(\mem[96] [0]), .B(data[0]), .S(n_97), .Z(n_106_80));
   MUX2_X1 i_106_0_720 (.A(\mem[97] [15]), .B(data[15]), .S(n_98), .Z(n_106_79));
   MUX2_X1 i_106_0_721 (.A(\mem[97] [14]), .B(data[14]), .S(n_98), .Z(n_106_78));
   MUX2_X1 i_106_0_722 (.A(\mem[97] [13]), .B(data[13]), .S(n_98), .Z(n_106_77));
   MUX2_X1 i_106_0_723 (.A(\mem[97] [12]), .B(data[12]), .S(n_98), .Z(n_106_76));
   MUX2_X1 i_106_0_724 (.A(\mem[97] [11]), .B(data[11]), .S(n_98), .Z(n_106_75));
   MUX2_X1 i_106_0_725 (.A(\mem[97] [10]), .B(data[10]), .S(n_98), .Z(n_106_74));
   MUX2_X1 i_106_0_726 (.A(\mem[97] [9]), .B(data[9]), .S(n_98), .Z(n_106_73));
   MUX2_X1 i_106_0_727 (.A(\mem[97] [8]), .B(data[8]), .S(n_98), .Z(n_106_72));
   MUX2_X1 i_106_0_728 (.A(\mem[97] [7]), .B(data[7]), .S(n_98), .Z(n_106_71));
   MUX2_X1 i_106_0_729 (.A(\mem[97] [6]), .B(data[6]), .S(n_98), .Z(n_106_70));
   MUX2_X1 i_106_0_730 (.A(\mem[97] [5]), .B(data[5]), .S(n_98), .Z(n_106_69));
   MUX2_X1 i_106_0_731 (.A(\mem[97] [4]), .B(data[4]), .S(n_98), .Z(n_106_68));
   MUX2_X1 i_106_0_732 (.A(\mem[97] [3]), .B(data[3]), .S(n_98), .Z(n_106_67));
   MUX2_X1 i_106_0_733 (.A(\mem[97] [2]), .B(data[2]), .S(n_98), .Z(n_106_66));
   MUX2_X1 i_106_0_734 (.A(\mem[97] [1]), .B(data[1]), .S(n_98), .Z(n_106_65));
   MUX2_X1 i_106_0_735 (.A(\mem[97] [0]), .B(data[0]), .S(n_98), .Z(n_106_64));
   MUX2_X1 i_106_0_736 (.A(\mem[98] [15]), .B(data[15]), .S(n_99), .Z(n_106_63));
   MUX2_X1 i_106_0_737 (.A(\mem[98] [14]), .B(data[14]), .S(n_99), .Z(n_106_62));
   MUX2_X1 i_106_0_738 (.A(\mem[98] [13]), .B(data[13]), .S(n_99), .Z(n_106_61));
   MUX2_X1 i_106_0_739 (.A(\mem[98] [12]), .B(data[12]), .S(n_99), .Z(n_106_60));
   MUX2_X1 i_106_0_740 (.A(\mem[98] [11]), .B(data[11]), .S(n_99), .Z(n_106_59));
   MUX2_X1 i_106_0_741 (.A(\mem[98] [10]), .B(data[10]), .S(n_99), .Z(n_106_58));
   MUX2_X1 i_106_0_742 (.A(\mem[98] [9]), .B(data[9]), .S(n_99), .Z(n_106_57));
   MUX2_X1 i_106_0_743 (.A(\mem[98] [8]), .B(data[8]), .S(n_99), .Z(n_106_56));
   MUX2_X1 i_106_0_744 (.A(\mem[98] [7]), .B(data[7]), .S(n_99), .Z(n_106_55));
   MUX2_X1 i_106_0_745 (.A(\mem[98] [6]), .B(data[6]), .S(n_99), .Z(n_106_54));
   MUX2_X1 i_106_0_746 (.A(\mem[98] [5]), .B(data[5]), .S(n_99), .Z(n_106_53));
   MUX2_X1 i_106_0_747 (.A(\mem[98] [4]), .B(data[4]), .S(n_99), .Z(n_106_52));
   MUX2_X1 i_106_0_748 (.A(\mem[98] [3]), .B(data[3]), .S(n_99), .Z(n_106_51));
   MUX2_X1 i_106_0_749 (.A(\mem[98] [2]), .B(data[2]), .S(n_99), .Z(n_106_50));
   MUX2_X1 i_106_0_750 (.A(\mem[98] [1]), .B(data[1]), .S(n_99), .Z(n_106_49));
   MUX2_X1 i_106_0_751 (.A(\mem[98] [0]), .B(data[0]), .S(n_99), .Z(n_106_48));
   MUX2_X1 i_106_0_752 (.A(\mem[99] [15]), .B(data[15]), .S(n_100), .Z(n_106_47));
   MUX2_X1 i_106_0_753 (.A(\mem[99] [14]), .B(data[14]), .S(n_100), .Z(n_106_46));
   MUX2_X1 i_106_0_754 (.A(\mem[99] [13]), .B(data[13]), .S(n_100), .Z(n_106_45));
   MUX2_X1 i_106_0_755 (.A(\mem[99] [12]), .B(data[12]), .S(n_100), .Z(n_106_44));
   MUX2_X1 i_106_0_756 (.A(\mem[99] [11]), .B(data[11]), .S(n_100), .Z(n_106_43));
   MUX2_X1 i_106_0_757 (.A(\mem[99] [10]), .B(data[10]), .S(n_100), .Z(n_106_42));
   MUX2_X1 i_106_0_758 (.A(\mem[99] [9]), .B(data[9]), .S(n_100), .Z(n_106_41));
   MUX2_X1 i_106_0_759 (.A(\mem[99] [8]), .B(data[8]), .S(n_100), .Z(n_106_40));
   MUX2_X1 i_106_0_760 (.A(\mem[99] [7]), .B(data[7]), .S(n_100), .Z(n_106_39));
   MUX2_X1 i_106_0_761 (.A(\mem[99] [6]), .B(data[6]), .S(n_100), .Z(n_106_38));
   MUX2_X1 i_106_0_762 (.A(\mem[99] [5]), .B(data[5]), .S(n_100), .Z(n_106_37));
   MUX2_X1 i_106_0_763 (.A(\mem[99] [4]), .B(data[4]), .S(n_100), .Z(n_106_36));
   MUX2_X1 i_106_0_764 (.A(\mem[99] [3]), .B(data[3]), .S(n_100), .Z(n_106_35));
   MUX2_X1 i_106_0_765 (.A(\mem[99] [2]), .B(data[2]), .S(n_100), .Z(n_106_34));
   MUX2_X1 i_106_0_766 (.A(\mem[99] [1]), .B(data[1]), .S(n_100), .Z(n_106_33));
   MUX2_X1 i_106_0_767 (.A(\mem[99] [0]), .B(data[0]), .S(n_100), .Z(n_106_32));
   MUX2_X1 i_106_0_768 (.A(\mem[100] [15]), .B(data[15]), .S(n_101), .Z(n_106_31));
   MUX2_X1 i_106_0_769 (.A(\mem[100] [14]), .B(data[14]), .S(n_101), .Z(n_106_30));
   MUX2_X1 i_106_0_770 (.A(\mem[100] [13]), .B(data[13]), .S(n_101), .Z(n_106_29));
   MUX2_X1 i_106_0_771 (.A(\mem[100] [12]), .B(data[12]), .S(n_101), .Z(n_106_28));
   MUX2_X1 i_106_0_772 (.A(\mem[100] [11]), .B(data[11]), .S(n_101), .Z(n_106_27));
   MUX2_X1 i_106_0_773 (.A(\mem[100] [10]), .B(data[10]), .S(n_101), .Z(n_106_26));
   MUX2_X1 i_106_0_774 (.A(\mem[100] [9]), .B(data[9]), .S(n_101), .Z(n_106_25));
   MUX2_X1 i_106_0_775 (.A(\mem[100] [8]), .B(data[8]), .S(n_101), .Z(n_106_24));
   MUX2_X1 i_106_0_776 (.A(\mem[100] [7]), .B(data[7]), .S(n_101), .Z(n_106_23));
   MUX2_X1 i_106_0_777 (.A(\mem[100] [6]), .B(data[6]), .S(n_101), .Z(n_106_22));
   MUX2_X1 i_106_0_778 (.A(\mem[100] [5]), .B(data[5]), .S(n_101), .Z(n_106_21));
   MUX2_X1 i_106_0_779 (.A(\mem[100] [4]), .B(data[4]), .S(n_101), .Z(n_106_20));
   MUX2_X1 i_106_0_780 (.A(\mem[100] [3]), .B(data[3]), .S(n_101), .Z(n_106_19));
   MUX2_X1 i_106_0_781 (.A(\mem[100] [2]), .B(data[2]), .S(n_101), .Z(n_106_18));
   MUX2_X1 i_106_0_782 (.A(\mem[100] [1]), .B(data[1]), .S(n_101), .Z(n_106_17));
   MUX2_X1 i_106_0_783 (.A(\mem[100] [0]), .B(data[0]), .S(n_101), .Z(n_106_16));
   MUX2_X1 i_106_0_784 (.A(\mem[0] [15]), .B(data[15]), .S(n_1), .Z(n_106_15));
   MUX2_X1 i_106_0_785 (.A(\mem[0] [14]), .B(data[14]), .S(n_1), .Z(n_106_14));
   MUX2_X1 i_106_0_786 (.A(\mem[0] [13]), .B(data[13]), .S(n_1), .Z(n_106_13));
   MUX2_X1 i_106_0_787 (.A(\mem[0] [12]), .B(data[12]), .S(n_1), .Z(n_106_12));
   MUX2_X1 i_106_0_788 (.A(\mem[0] [11]), .B(data[11]), .S(n_1), .Z(n_106_11));
   MUX2_X1 i_106_0_789 (.A(\mem[0] [10]), .B(data[10]), .S(n_1), .Z(n_106_10));
   MUX2_X1 i_106_0_790 (.A(\mem[0] [9]), .B(data[9]), .S(n_1), .Z(n_106_9));
   MUX2_X1 i_106_0_791 (.A(\mem[0] [8]), .B(data[8]), .S(n_1), .Z(n_106_8));
   MUX2_X1 i_106_0_792 (.A(\mem[0] [7]), .B(data[7]), .S(n_1), .Z(n_106_7));
   MUX2_X1 i_106_0_793 (.A(\mem[0] [6]), .B(data[6]), .S(n_1), .Z(n_106_6));
   MUX2_X1 i_106_0_794 (.A(\mem[0] [5]), .B(data[5]), .S(n_1), .Z(n_106_5));
   MUX2_X1 i_106_0_795 (.A(\mem[0] [4]), .B(data[4]), .S(n_1), .Z(n_106_4));
   MUX2_X1 i_106_0_796 (.A(\mem[0] [3]), .B(data[3]), .S(n_1), .Z(n_106_3));
   MUX2_X1 i_106_0_797 (.A(\mem[0] [2]), .B(data[2]), .S(n_1), .Z(n_106_2));
   MUX2_X1 i_106_0_798 (.A(\mem[0] [1]), .B(data[1]), .S(n_1), .Z(n_106_1));
   MUX2_X1 i_106_0_799 (.A(\mem[0] [0]), .B(data[0]), .S(n_1), .Z(n_106_0));
   DFF_X1 \temp_reg[15]  (.D(n_1_15), .CK(n_0), .Q(dataout[15]), .QN());
   DFF_X1 \temp_reg[14]  (.D(n_1_14), .CK(n_0), .Q(dataout[14]), .QN());
   DFF_X1 \temp_reg[13]  (.D(n_1_13), .CK(n_0), .Q(dataout[13]), .QN());
   DFF_X1 \temp_reg[12]  (.D(n_1_12), .CK(n_0), .Q(dataout[12]), .QN());
   DFF_X1 \temp_reg[11]  (.D(n_1_11), .CK(n_0), .Q(dataout[11]), .QN());
   DFF_X1 \temp_reg[10]  (.D(n_1_10), .CK(n_0), .Q(dataout[10]), .QN());
   DFF_X1 \temp_reg[9]  (.D(n_1_9), .CK(n_0), .Q(dataout[9]), .QN());
   DFF_X1 \temp_reg[8]  (.D(n_1_8), .CK(n_0), .Q(dataout[8]), .QN());
   DFF_X1 \temp_reg[7]  (.D(n_1_7), .CK(n_0), .Q(dataout[7]), .QN());
   DFF_X1 \temp_reg[6]  (.D(n_1_6), .CK(n_0), .Q(dataout[6]), .QN());
   DFF_X1 \temp_reg[5]  (.D(n_1_5), .CK(n_0), .Q(dataout[5]), .QN());
   DFF_X1 \temp_reg[4]  (.D(n_1_4), .CK(n_0), .Q(dataout[4]), .QN());
   DFF_X1 \temp_reg[3]  (.D(n_1_3), .CK(n_0), .Q(dataout[3]), .QN());
   DFF_X1 \temp_reg[2]  (.D(n_1_2), .CK(n_0), .Q(dataout[2]), .QN());
   DFF_X1 \temp_reg[1]  (.D(n_1_1), .CK(n_0), .Q(dataout[1]), .QN());
   DFF_X1 \temp_reg[0]  (.D(n_1_0), .CK(n_0), .Q(dataout[0]), .QN());
   INV_X1 i_1_0_0 (.A(clk), .ZN(n_0));
   MUX2_X1 i_1_1_0 (.A(dataout[0]), .B(n_1_1_0), .S(read_signal), .Z(n_1_0));
   NAND4_X1 i_1_1_1 (.A1(n_1_1_14), .A2(n_1_1_12), .A3(n_1_1_7), .A4(n_1_1_1), 
      .ZN(n_1_1_0));
   AOI221_X1 i_1_1_2 (.A(n_1_1_2), .B1(n_1_1_1052), .B2(\mem[23] [0]), .C1(
      \mem[87] [0]), .C2(n_1_1_1144), .ZN(n_1_1_1));
   NAND4_X1 i_1_1_3 (.A1(n_1_1_49), .A2(n_1_1_40), .A3(n_1_1_4), .A4(n_1_1_3), 
      .ZN(n_1_1_2));
   AOI222_X1 i_1_1_4 (.A1(\mem[61] [0]), .A2(n_1_1_1057), .B1(n_1_1_1046), 
      .B2(\mem[60] [0]), .C1(\mem[13] [0]), .C2(n_1_1_1075), .ZN(n_1_1_3));
   AOI221_X1 i_1_1_5 (.A(n_1_1_5), .B1(n_1_1_1088), .B2(\mem[31] [0]), .C1(
      \mem[71] [0]), .C2(n_1_1_1126), .ZN(n_1_1_4));
   NAND3_X1 i_1_1_6 (.A1(n_1_1_42), .A2(n_1_1_41), .A3(n_1_1_6), .ZN(n_1_1_5));
   AOI22_X1 i_1_1_7 (.A1(\mem[72] [0]), .A2(n_1_1_1127), .B1(n_1_1_1074), 
      .B2(\mem[9] [0]), .ZN(n_1_1_6));
   NOR4_X1 i_1_1_8 (.A1(n_1_1_11), .A2(n_1_1_10), .A3(n_1_1_9), .A4(n_1_1_8), 
      .ZN(n_1_1_7));
   NAND4_X1 i_1_1_9 (.A1(n_1_1_64), .A2(n_1_1_58), .A3(n_1_1_57), .A4(n_1_1_36), 
      .ZN(n_1_1_8));
   NAND4_X1 i_1_1_10 (.A1(n_1_1_65), .A2(n_1_1_50), .A3(n_1_1_35), .A4(n_1_1_33), 
      .ZN(n_1_1_9));
   NAND4_X1 i_1_1_11 (.A1(n_1_1_55), .A2(n_1_1_51), .A3(n_1_1_38), .A4(n_1_1_37), 
      .ZN(n_1_1_10));
   NAND4_X1 i_1_1_12 (.A1(n_1_1_61), .A2(n_1_1_56), .A3(n_1_1_54), .A4(n_1_1_34), 
      .ZN(n_1_1_11));
   AOI221_X1 i_1_1_13 (.A(n_1_1_13), .B1(n_1_1_1031), .B2(\mem[39] [0]), 
      .C1(\mem[75] [0]), .C2(n_1_1_1061), .ZN(n_1_1_12));
   NAND3_X1 i_1_1_14 (.A1(n_1_1_46), .A2(n_1_1_29), .A3(n_1_1_28), .ZN(n_1_1_13));
   AOI221_X1 i_1_1_15 (.A(n_1_1_15), .B1(n_1_1_1035), .B2(\mem[50] [0]), 
      .C1(\mem[86] [0]), .C2(n_1_1_1142), .ZN(n_1_1_14));
   NAND3_X1 i_1_1_16 (.A1(n_1_1_47), .A2(n_1_1_18), .A3(n_1_1_16), .ZN(n_1_1_15));
   AOI221_X1 i_1_1_17 (.A(n_1_1_17), .B1(n_1_1_1070), .B2(\mem[4] [0]), .C1(
      \mem[55] [0]), .C2(n_1_1_1107), .ZN(n_1_1_16));
   NAND3_X1 i_1_1_18 (.A1(n_1_1_62), .A2(n_1_1_30), .A3(n_1_1_24), .ZN(n_1_1_17));
   NOR4_X1 i_1_1_19 (.A1(n_1_1_22), .A2(n_1_1_21), .A3(n_1_1_20), .A4(n_1_1_19), 
      .ZN(n_1_1_18));
   NAND4_X1 i_1_1_20 (.A1(n_1_1_48), .A2(n_1_1_27), .A3(n_1_1_26), .A4(n_1_1_25), 
      .ZN(n_1_1_19));
   NAND4_X1 i_1_1_21 (.A1(n_1_1_63), .A2(n_1_1_52), .A3(n_1_1_44), .A4(n_1_1_31), 
      .ZN(n_1_1_20));
   NAND4_X1 i_1_1_22 (.A1(n_1_1_60), .A2(n_1_1_59), .A3(n_1_1_45), .A4(n_1_1_32), 
      .ZN(n_1_1_21));
   NAND4_X1 i_1_1_23 (.A1(n_1_1_53), .A2(n_1_1_43), .A3(n_1_1_39), .A4(n_1_1_23), 
      .ZN(n_1_1_22));
   AOI22_X1 i_1_1_24 (.A1(\mem[54] [0]), .A2(n_1_1_1106), .B1(n_1_1_1030), 
      .B2(\mem[20] [0]), .ZN(n_1_1_23));
   AOI22_X1 i_1_1_25 (.A1(\mem[66] [0]), .A2(n_1_1_1120), .B1(n_1_1_1064), 
      .B2(\mem[18] [0]), .ZN(n_1_1_24));
   AOI22_X1 i_1_1_26 (.A1(\mem[79] [0]), .A2(n_1_1_1135), .B1(n_1_1_1050), 
      .B2(\mem[90] [0]), .ZN(n_1_1_25));
   AOI22_X1 i_1_1_27 (.A1(\mem[65] [0]), .A2(n_1_1_1119), .B1(n_1_1_1109), 
      .B2(\mem[58] [0]), .ZN(n_1_1_26));
   AOI22_X1 i_1_1_28 (.A1(\mem[93] [0]), .A2(n_1_1_1155), .B1(n_1_1_1039), 
      .B2(\mem[76] [0]), .ZN(n_1_1_27));
   AOI22_X1 i_1_1_29 (.A1(\mem[41] [0]), .A2(n_1_1_1100), .B1(n_1_1_1096), 
      .B2(\mem[37] [0]), .ZN(n_1_1_28));
   AOI22_X1 i_1_1_30 (.A1(\mem[57] [0]), .A2(n_1_1_1108), .B1(n_1_1_1048), 
      .B2(\mem[10] [0]), .ZN(n_1_1_29));
   AOI22_X1 i_1_1_31 (.A1(\mem[48] [0]), .A2(n_1_1_1104), .B1(n_1_1_1087), 
      .B2(\mem[30] [0]), .ZN(n_1_1_30));
   AOI22_X1 i_1_1_32 (.A1(\mem[100] [0]), .A2(n_1_1_1174), .B1(n_1_1_1038), 
      .B2(\mem[15] [0]), .ZN(n_1_1_31));
   AOI22_X1 i_1_1_33 (.A1(\mem[94] [0]), .A2(n_1_1_1157), .B1(n_1_1_1041), 
      .B2(\mem[7] [0]), .ZN(n_1_1_32));
   AOI22_X1 i_1_1_34 (.A1(\mem[40] [0]), .A2(n_1_1_1099), .B1(n_1_1_1058), 
      .B2(\mem[85] [0]), .ZN(n_1_1_33));
   AOI22_X1 i_1_1_35 (.A1(\mem[70] [0]), .A2(n_1_1_1125), .B1(n_1_1_1123), 
      .B2(\mem[69] [0]), .ZN(n_1_1_34));
   AOI22_X1 i_1_1_36 (.A1(\mem[5] [0]), .A2(n_1_1_1071), .B1(n_1_1_1063), 
      .B2(\mem[11] [0]), .ZN(n_1_1_35));
   AOI22_X1 i_1_1_37 (.A1(\mem[32] [0]), .A2(n_1_1_1091), .B1(n_1_1_1043), 
      .B2(\mem[53] [0]), .ZN(n_1_1_36));
   AOI22_X1 i_1_1_38 (.A1(\mem[96] [0]), .A2(n_1_1_1163), .B1(n_1_1_1051), 
      .B2(\mem[29] [0]), .ZN(n_1_1_37));
   AOI22_X1 i_1_1_39 (.A1(\mem[92] [0]), .A2(n_1_1_1153), .B1(n_1_1_1111), 
      .B2(\mem[59] [0]), .ZN(n_1_1_38));
   AOI22_X1 i_1_1_40 (.A1(\mem[84] [0]), .A2(n_1_1_1062), .B1(n_1_1_1028), 
      .B2(\mem[82] [0]), .ZN(n_1_1_39));
   AOI22_X1 i_1_1_41 (.A1(\mem[68] [0]), .A2(n_1_1_1122), .B1(n_1_1_1044), 
      .B2(\mem[26] [0]), .ZN(n_1_1_40));
   AOI22_X1 i_1_1_42 (.A1(\mem[35] [0]), .A2(n_1_1_1094), .B1(n_1_1_1073), 
      .B2(\mem[8] [0]), .ZN(n_1_1_41));
   AOI22_X1 i_1_1_43 (.A1(\mem[88] [0]), .A2(n_1_1_1056), .B1(n_1_1_1036), 
      .B2(\mem[14] [0]), .ZN(n_1_1_42));
   AOI22_X1 i_1_1_44 (.A1(\mem[21] [0]), .A2(n_1_1_1081), .B1(n_1_1_1069), 
      .B2(\mem[3] [0]), .ZN(n_1_1_43));
   AOI22_X1 i_1_1_45 (.A1(\mem[25] [0]), .A2(n_1_1_1084), .B1(n_1_1_1078), 
      .B2(\mem[16] [0]), .ZN(n_1_1_44));
   AOI22_X1 i_1_1_46 (.A1(\mem[33] [0]), .A2(n_1_1_1092), .B1(n_1_1_1080), 
      .B2(\mem[19] [0]), .ZN(n_1_1_45));
   AOI22_X1 i_1_1_47 (.A1(\mem[73] [0]), .A2(n_1_1_1129), .B1(n_1_1_1101), 
      .B2(\mem[46] [0]), .ZN(n_1_1_46));
   AOI22_X1 i_1_1_48 (.A1(\mem[52] [0]), .A2(n_1_1_1040), .B1(n_1_1_1025), 
      .B2(\mem[43] [0]), .ZN(n_1_1_47));
   AOI22_X1 i_1_1_49 (.A1(\mem[78] [0]), .A2(n_1_1_1134), .B1(n_1_1_1068), 
      .B2(\mem[2] [0]), .ZN(n_1_1_48));
   AOI22_X1 i_1_1_50 (.A1(\mem[49] [0]), .A2(n_1_1_1105), .B1(n_1_1_1055), 
      .B2(\mem[74] [0]), .ZN(n_1_1_49));
   AOI22_X1 i_1_1_51 (.A1(\mem[97] [0]), .A2(n_1_1_1165), .B1(n_1_1_1093), 
      .B2(\mem[34] [0]), .ZN(n_1_1_50));
   AOI22_X1 i_1_1_52 (.A1(\mem[47] [0]), .A2(n_1_1_1102), .B1(n_1_1_1026), 
      .B2(\mem[56] [0]), .ZN(n_1_1_51));
   AOI22_X1 i_1_1_53 (.A1(\mem[38] [0]), .A2(n_1_1_1097), .B1(n_1_1_1033), 
      .B2(\mem[42] [0]), .ZN(n_1_1_52));
   AOI22_X1 i_1_1_54 (.A1(\mem[51] [0]), .A2(n_1_1_1059), .B1(n_1_1_1054), 
      .B2(\mem[22] [0]), .ZN(n_1_1_53));
   AOI22_X1 i_1_1_55 (.A1(\mem[89] [0]), .A2(n_1_1_1148), .B1(n_1_1_1121), 
      .B2(\mem[67] [0]), .ZN(n_1_1_54));
   AOI22_X1 i_1_1_56 (.A1(\mem[95] [0]), .A2(n_1_1_1053), .B1(n_1_1_1047), 
      .B2(\mem[83] [0]), .ZN(n_1_1_55));
   AOI22_X1 i_1_1_57 (.A1(\mem[77] [0]), .A2(n_1_1_1133), .B1(n_1_1_1072), 
      .B2(\mem[6] [0]), .ZN(n_1_1_56));
   AOI22_X1 i_1_1_58 (.A1(\mem[36] [0]), .A2(n_1_1_1095), .B1(n_1_1_1049), 
      .B2(\mem[17] [0]), .ZN(n_1_1_57));
   AOI22_X1 i_1_1_59 (.A1(\mem[80] [0]), .A2(n_1_1_1138), .B1(n_1_1_1042), 
      .B2(\mem[12] [0]), .ZN(n_1_1_58));
   AOI22_X1 i_1_1_60 (.A1(\mem[99] [0]), .A2(n_1_1_1171), .B1(n_1_1_1066), 
      .B2(\mem[0] [0]), .ZN(n_1_1_59));
   AOI22_X1 i_1_1_61 (.A1(\mem[81] [0]), .A2(n_1_1_1139), .B1(n_1_1_1027), 
      .B2(\mem[27] [0]), .ZN(n_1_1_60));
   AOI22_X1 i_1_1_62 (.A1(\mem[98] [0]), .A2(n_1_1_1168), .B1(n_1_1_1060), 
      .B2(\mem[28] [0]), .ZN(n_1_1_61));
   AOI22_X1 i_1_1_63 (.A1(\mem[64] [0]), .A2(n_1_1_1118), .B1(n_1_1_1032), 
      .B2(\mem[44] [0]), .ZN(n_1_1_62));
   AOI22_X1 i_1_1_64 (.A1(\mem[45] [0]), .A2(n_1_1_1045), .B1(n_1_1_1037), 
      .B2(\mem[91] [0]), .ZN(n_1_1_63));
   AOI22_X1 i_1_1_65 (.A1(\mem[63] [0]), .A2(n_1_1_1116), .B1(n_1_1_1083), 
      .B2(\mem[24] [0]), .ZN(n_1_1_64));
   AOI22_X1 i_1_1_66 (.A1(\mem[1] [0]), .A2(n_1_1_1067), .B1(n_1_1_1029), 
      .B2(\mem[62] [0]), .ZN(n_1_1_65));
   INV_X1 i_1_1_67 (.A(n_1_1_66), .ZN(n_1_1));
   OAI22_X1 i_1_1_68 (.A1(n_1_1_103), .A2(n_1_1_67), .B1(read_signal), .B2(
      dataout[1]), .ZN(n_1_1_66));
   NAND4_X1 i_1_1_69 (.A1(n_1_1_102), .A2(n_1_1_88), .A3(n_1_1_83), .A4(n_1_1_68), 
      .ZN(n_1_1_67));
   NOR4_X1 i_1_1_70 (.A1(n_1_1_78), .A2(n_1_1_74), .A3(n_1_1_72), .A4(n_1_1_69), 
      .ZN(n_1_1_68));
   NAND4_X1 i_1_1_71 (.A1(n_1_1_128), .A2(n_1_1_127), .A3(n_1_1_71), .A4(
      n_1_1_70), .ZN(n_1_1_69));
   AOI22_X1 i_1_1_72 (.A1(\mem[81] [1]), .A2(n_1_1_1139), .B1(n_1_1_1104), 
      .B2(\mem[48] [1]), .ZN(n_1_1_70));
   AOI22_X1 i_1_1_73 (.A1(\mem[75] [1]), .A2(n_1_1_1061), .B1(n_1_1_1048), 
      .B2(\mem[10] [1]), .ZN(n_1_1_71));
   NAND3_X1 i_1_1_74 (.A1(read_signal), .A2(n_1_1_126), .A3(n_1_1_73), .ZN(
      n_1_1_72));
   AOI222_X1 i_1_1_75 (.A1(\mem[96] [1]), .A2(n_1_1_1163), .B1(n_1_1_1081), 
      .B2(\mem[21] [1]), .C1(n_1_1_1051), .C2(\mem[29] [1]), .ZN(n_1_1_73));
   NAND4_X1 i_1_1_76 (.A1(n_1_1_130), .A2(n_1_1_77), .A3(n_1_1_76), .A4(n_1_1_75), 
      .ZN(n_1_1_74));
   AOI22_X1 i_1_1_77 (.A1(\mem[85] [1]), .A2(n_1_1_1058), .B1(n_1_1_1036), 
      .B2(\mem[14] [1]), .ZN(n_1_1_75));
   AOI22_X1 i_1_1_78 (.A1(\mem[2] [1]), .A2(n_1_1_1068), .B1(n_1_1_1050), 
      .B2(\mem[90] [1]), .ZN(n_1_1_76));
   AOI22_X1 i_1_1_79 (.A1(\mem[94] [1]), .A2(n_1_1_1157), .B1(n_1_1_1105), 
      .B2(\mem[49] [1]), .ZN(n_1_1_77));
   NAND4_X1 i_1_1_80 (.A1(n_1_1_82), .A2(n_1_1_81), .A3(n_1_1_80), .A4(n_1_1_79), 
      .ZN(n_1_1_78));
   AOI22_X1 i_1_1_81 (.A1(\mem[80] [1]), .A2(n_1_1_1138), .B1(n_1_1_1119), 
      .B2(\mem[65] [1]), .ZN(n_1_1_79));
   AOI22_X1 i_1_1_82 (.A1(\mem[66] [1]), .A2(n_1_1_1120), .B1(n_1_1_1026), 
      .B2(\mem[56] [1]), .ZN(n_1_1_80));
   AOI22_X1 i_1_1_83 (.A1(\mem[12] [1]), .A2(n_1_1_1042), .B1(n_1_1_1032), 
      .B2(\mem[44] [1]), .ZN(n_1_1_81));
   AOI22_X1 i_1_1_84 (.A1(\mem[63] [1]), .A2(n_1_1_1116), .B1(n_1_1_1071), 
      .B2(\mem[5] [1]), .ZN(n_1_1_82));
   AOI221_X1 i_1_1_85 (.A(n_1_1_84), .B1(n_1_1_1165), .B2(\mem[97] [1]), 
      .C1(\mem[99] [1]), .C2(n_1_1_1171), .ZN(n_1_1_83));
   NAND3_X1 i_1_1_86 (.A1(n_1_1_87), .A2(n_1_1_86), .A3(n_1_1_85), .ZN(n_1_1_84));
   AOI22_X1 i_1_1_87 (.A1(\mem[59] [1]), .A2(n_1_1_1111), .B1(n_1_1_1046), 
      .B2(\mem[60] [1]), .ZN(n_1_1_85));
   AOI22_X1 i_1_1_88 (.A1(\mem[79] [1]), .A2(n_1_1_1135), .B1(n_1_1_1044), 
      .B2(\mem[26] [1]), .ZN(n_1_1_86));
   AOI22_X1 i_1_1_89 (.A1(\mem[47] [1]), .A2(n_1_1_1102), .B1(n_1_1_1083), 
      .B2(\mem[24] [1]), .ZN(n_1_1_87));
   AOI221_X1 i_1_1_90 (.A(n_1_1_89), .B1(n_1_1_1063), .B2(\mem[11] [1]), 
      .C1(\mem[64] [1]), .C2(n_1_1_1118), .ZN(n_1_1_88));
   NAND4_X1 i_1_1_91 (.A1(n_1_1_98), .A2(n_1_1_94), .A3(n_1_1_91), .A4(n_1_1_90), 
      .ZN(n_1_1_89));
   AOI222_X1 i_1_1_92 (.A1(\mem[86] [1]), .A2(n_1_1_1142), .B1(n_1_1_1091), 
      .B2(\mem[32] [1]), .C1(n_1_1_1060), .C2(\mem[28] [1]), .ZN(n_1_1_90));
   AOI221_X1 i_1_1_93 (.A(n_1_1_92), .B1(n_1_1_1033), .B2(\mem[42] [1]), 
      .C1(\mem[58] [1]), .C2(n_1_1_1109), .ZN(n_1_1_91));
   NAND3_X1 i_1_1_94 (.A1(n_1_1_129), .A2(n_1_1_125), .A3(n_1_1_93), .ZN(
      n_1_1_92));
   AOI22_X1 i_1_1_95 (.A1(\mem[40] [1]), .A2(n_1_1_1099), .B1(n_1_1_1062), 
      .B2(\mem[84] [1]), .ZN(n_1_1_93));
   AOI221_X1 i_1_1_96 (.A(n_1_1_95), .B1(n_1_1_1031), .B2(\mem[39] [1]), 
      .C1(\mem[51] [1]), .C2(n_1_1_1059), .ZN(n_1_1_94));
   NAND2_X1 i_1_1_97 (.A1(n_1_1_97), .A2(n_1_1_96), .ZN(n_1_1_95));
   AOI222_X1 i_1_1_98 (.A1(\mem[83] [1]), .A2(n_1_1_1047), .B1(n_1_1_1025), 
      .B2(\mem[43] [1]), .C1(\mem[30] [1]), .C2(n_1_1_1087), .ZN(n_1_1_96));
   AOI222_X1 i_1_1_99 (.A1(\mem[98] [1]), .A2(n_1_1_1168), .B1(n_1_1_1125), 
      .B2(\mem[70] [1]), .C1(n_1_1_1094), .C2(\mem[35] [1]), .ZN(n_1_1_97));
   AOI221_X1 i_1_1_100 (.A(n_1_1_99), .B1(n_1_1_1080), .B2(\mem[19] [1]), 
      .C1(\mem[45] [1]), .C2(n_1_1_1045), .ZN(n_1_1_98));
   NAND3_X1 i_1_1_101 (.A1(n_1_1_124), .A2(n_1_1_101), .A3(n_1_1_100), .ZN(
      n_1_1_99));
   AOI22_X1 i_1_1_102 (.A1(\mem[16] [1]), .A2(n_1_1_1078), .B1(n_1_1_1064), 
      .B2(\mem[18] [1]), .ZN(n_1_1_100));
   AOI22_X1 i_1_1_103 (.A1(\mem[25] [1]), .A2(n_1_1_1084), .B1(n_1_1_1052), 
      .B2(\mem[23] [1]), .ZN(n_1_1_101));
   AOI222_X1 i_1_1_104 (.A1(\mem[93] [1]), .A2(n_1_1_1155), .B1(n_1_1_1134), 
      .B2(\mem[78] [1]), .C1(n_1_1_1073), .C2(\mem[8] [1]), .ZN(n_1_1_102));
   NAND4_X1 i_1_1_105 (.A1(n_1_1_119), .A2(n_1_1_114), .A3(n_1_1_109), .A4(
      n_1_1_104), .ZN(n_1_1_103));
   AOI221_X1 i_1_1_106 (.A(n_1_1_105), .B1(n_1_1_1092), .B2(\mem[33] [1]), 
      .C1(\mem[74] [1]), .C2(n_1_1_1055), .ZN(n_1_1_104));
   NAND3_X1 i_1_1_107 (.A1(n_1_1_108), .A2(n_1_1_107), .A3(n_1_1_106), .ZN(
      n_1_1_105));
   AOI22_X1 i_1_1_108 (.A1(\mem[72] [1]), .A2(n_1_1_1127), .B1(n_1_1_1028), 
      .B2(\mem[82] [1]), .ZN(n_1_1_106));
   AOI22_X1 i_1_1_109 (.A1(\mem[37] [1]), .A2(n_1_1_1096), .B1(n_1_1_1057), 
      .B2(\mem[61] [1]), .ZN(n_1_1_107));
   AOI22_X1 i_1_1_110 (.A1(\mem[4] [1]), .A2(n_1_1_1070), .B1(n_1_1_1030), 
      .B2(\mem[20] [1]), .ZN(n_1_1_108));
   AOI221_X1 i_1_1_111 (.A(n_1_1_110), .B1(n_1_1_1069), .B2(\mem[3] [1]), 
      .C1(\mem[89] [1]), .C2(n_1_1_1148), .ZN(n_1_1_109));
   NAND3_X1 i_1_1_112 (.A1(n_1_1_113), .A2(n_1_1_112), .A3(n_1_1_111), .ZN(
      n_1_1_110));
   AOI22_X1 i_1_1_113 (.A1(\mem[71] [1]), .A2(n_1_1_1126), .B1(n_1_1_1107), 
      .B2(\mem[55] [1]), .ZN(n_1_1_111));
   AOI22_X1 i_1_1_114 (.A1(\mem[67] [1]), .A2(n_1_1_1121), .B1(n_1_1_1049), 
      .B2(\mem[17] [1]), .ZN(n_1_1_112));
   AOI22_X1 i_1_1_115 (.A1(\mem[87] [1]), .A2(n_1_1_1144), .B1(n_1_1_1100), 
      .B2(\mem[41] [1]), .ZN(n_1_1_113));
   AOI221_X1 i_1_1_116 (.A(n_1_1_115), .B1(n_1_1_1093), .B2(\mem[34] [1]), 
      .C1(\mem[46] [1]), .C2(n_1_1_1101), .ZN(n_1_1_114));
   NAND3_X1 i_1_1_117 (.A1(n_1_1_118), .A2(n_1_1_117), .A3(n_1_1_116), .ZN(
      n_1_1_115));
   AOI22_X1 i_1_1_118 (.A1(\mem[91] [1]), .A2(n_1_1_1037), .B1(n_1_1_1035), 
      .B2(\mem[50] [1]), .ZN(n_1_1_116));
   AOI22_X1 i_1_1_119 (.A1(\mem[100] [1]), .A2(n_1_1_1174), .B1(n_1_1_1054), 
      .B2(\mem[22] [1]), .ZN(n_1_1_117));
   AOI22_X1 i_1_1_120 (.A1(\mem[69] [1]), .A2(n_1_1_1123), .B1(n_1_1_1041), 
      .B2(\mem[7] [1]), .ZN(n_1_1_118));
   AOI221_X1 i_1_1_121 (.A(n_1_1_120), .B1(n_1_1_1067), .B2(\mem[1] [1]), 
      .C1(\mem[38] [1]), .C2(n_1_1_1097), .ZN(n_1_1_119));
   NAND3_X1 i_1_1_122 (.A1(n_1_1_123), .A2(n_1_1_122), .A3(n_1_1_121), .ZN(
      n_1_1_120));
   AOI22_X1 i_1_1_123 (.A1(\mem[77] [1]), .A2(n_1_1_1133), .B1(n_1_1_1038), 
      .B2(\mem[15] [1]), .ZN(n_1_1_121));
   AOI22_X1 i_1_1_124 (.A1(\mem[92] [1]), .A2(n_1_1_1153), .B1(n_1_1_1095), 
      .B2(\mem[36] [1]), .ZN(n_1_1_122));
   AOI22_X1 i_1_1_125 (.A1(\mem[73] [1]), .A2(n_1_1_1129), .B1(n_1_1_1074), 
      .B2(\mem[9] [1]), .ZN(n_1_1_123));
   AOI22_X1 i_1_1_126 (.A1(\mem[6] [1]), .A2(n_1_1_1072), .B1(n_1_1_1053), 
      .B2(\mem[95] [1]), .ZN(n_1_1_124));
   AOI22_X1 i_1_1_127 (.A1(\mem[53] [1]), .A2(n_1_1_1043), .B1(n_1_1_1039), 
      .B2(\mem[76] [1]), .ZN(n_1_1_125));
   AOI22_X1 i_1_1_128 (.A1(\mem[57] [1]), .A2(n_1_1_1108), .B1(n_1_1_1106), 
      .B2(\mem[54] [1]), .ZN(n_1_1_126));
   AOI22_X1 i_1_1_129 (.A1(\mem[68] [1]), .A2(n_1_1_1122), .B1(n_1_1_1075), 
      .B2(\mem[13] [1]), .ZN(n_1_1_127));
   AOI22_X1 i_1_1_130 (.A1(\mem[0] [1]), .A2(n_1_1_1066), .B1(n_1_1_1040), 
      .B2(\mem[52] [1]), .ZN(n_1_1_128));
   AOI22_X1 i_1_1_131 (.A1(\mem[88] [1]), .A2(n_1_1_1056), .B1(n_1_1_1029), 
      .B2(\mem[62] [1]), .ZN(n_1_1_129));
   AOI22_X1 i_1_1_132 (.A1(\mem[31] [1]), .A2(n_1_1_1088), .B1(n_1_1_1027), 
      .B2(\mem[27] [1]), .ZN(n_1_1_130));
   AOI21_X1 i_1_1_133 (.A(n_1_1_192), .B1(n_1_1_131), .B2(read_signal), .ZN(
      n_1_2));
   AOI221_X1 i_1_1_134 (.A(n_1_1_132), .B1(n_1_1_1045), .B2(\mem[45] [2]), 
      .C1(\mem[89] [2]), .C2(n_1_1_1148), .ZN(n_1_1_131));
   NAND4_X1 i_1_1_135 (.A1(n_1_1_164), .A2(n_1_1_143), .A3(n_1_1_139), .A4(
      n_1_1_133), .ZN(n_1_1_132));
   AOI221_X1 i_1_1_136 (.A(n_1_1_134), .B1(n_1_1_1066), .B2(\mem[0] [2]), 
      .C1(\mem[66] [2]), .C2(n_1_1_1120), .ZN(n_1_1_133));
   NAND3_X1 i_1_1_137 (.A1(n_1_1_138), .A2(n_1_1_137), .A3(n_1_1_135), .ZN(
      n_1_1_134));
   AOI221_X1 i_1_1_138 (.A(n_1_1_136), .B1(n_1_1_1101), .B2(\mem[46] [2]), 
      .C1(\mem[72] [2]), .C2(n_1_1_1127), .ZN(n_1_1_135));
   NAND3_X1 i_1_1_139 (.A1(n_1_1_180), .A2(n_1_1_179), .A3(n_1_1_178), .ZN(
      n_1_1_136));
   AOI22_X1 i_1_1_140 (.A1(\mem[32] [2]), .A2(n_1_1_1091), .B1(n_1_1_1075), 
      .B2(\mem[13] [2]), .ZN(n_1_1_137));
   AOI222_X1 i_1_1_141 (.A1(\mem[68] [2]), .A2(n_1_1_1122), .B1(n_1_1_1095), 
      .B2(\mem[36] [2]), .C1(n_1_1_1057), .C2(\mem[61] [2]), .ZN(n_1_1_138));
   AOI221_X1 i_1_1_142 (.A(n_1_1_140), .B1(n_1_1_1064), .B2(\mem[18] [2]), 
      .C1(\mem[74] [2]), .C2(n_1_1_1055), .ZN(n_1_1_139));
   NAND4_X1 i_1_1_143 (.A1(n_1_1_176), .A2(n_1_1_175), .A3(n_1_1_142), .A4(
      n_1_1_141), .ZN(n_1_1_140));
   AOI222_X1 i_1_1_144 (.A1(\mem[73] [2]), .A2(n_1_1_1129), .B1(n_1_1_1111), 
      .B2(\mem[59] [2]), .C1(n_1_1_1048), .C2(\mem[10] [2]), .ZN(n_1_1_141));
   AOI22_X1 i_1_1_145 (.A1(\mem[86] [2]), .A2(n_1_1_1142), .B1(n_1_1_1032), 
      .B2(\mem[44] [2]), .ZN(n_1_1_142));
   AOI221_X1 i_1_1_146 (.A(n_1_1_144), .B1(n_1_1_1059), .B2(\mem[51] [2]), 
      .C1(\mem[57] [2]), .C2(n_1_1_1108), .ZN(n_1_1_143));
   NAND4_X1 i_1_1_147 (.A1(n_1_1_185), .A2(n_1_1_163), .A3(n_1_1_161), .A4(
      n_1_1_145), .ZN(n_1_1_144));
   NOR4_X1 i_1_1_148 (.A1(n_1_1_158), .A2(n_1_1_149), .A3(n_1_1_148), .A4(
      n_1_1_146), .ZN(n_1_1_145));
   NAND4_X1 i_1_1_149 (.A1(n_1_1_187), .A2(n_1_1_184), .A3(n_1_1_177), .A4(
      n_1_1_147), .ZN(n_1_1_146));
   AOI22_X1 i_1_1_150 (.A1(\mem[28] [2]), .A2(n_1_1_1060), .B1(n_1_1_1050), 
      .B2(\mem[90] [2]), .ZN(n_1_1_147));
   NAND4_X1 i_1_1_151 (.A1(n_1_1_191), .A2(n_1_1_183), .A3(n_1_1_181), .A4(
      n_1_1_169), .ZN(n_1_1_148));
   NAND4_X1 i_1_1_152 (.A1(n_1_1_155), .A2(n_1_1_152), .A3(n_1_1_151), .A4(
      n_1_1_150), .ZN(n_1_1_149));
   AOI222_X1 i_1_1_153 (.A1(\mem[63] [2]), .A2(n_1_1_1116), .B1(n_1_1_1087), 
      .B2(\mem[30] [2]), .C1(n_1_1_1037), .C2(\mem[91] [2]), .ZN(n_1_1_150));
   AOI222_X1 i_1_1_154 (.A1(\mem[65] [2]), .A2(n_1_1_1119), .B1(n_1_1_1052), 
      .B2(\mem[23] [2]), .C1(n_1_1_1049), .C2(\mem[17] [2]), .ZN(n_1_1_151));
   AOI221_X1 i_1_1_155 (.A(n_1_1_153), .B1(n_1_1_1042), .B2(\mem[12] [2]), 
      .C1(\mem[47] [2]), .C2(n_1_1_1102), .ZN(n_1_1_152));
   NAND4_X1 i_1_1_156 (.A1(n_1_1_170), .A2(n_1_1_166), .A3(n_1_1_165), .A4(
      n_1_1_154), .ZN(n_1_1_153));
   AOI22_X1 i_1_1_157 (.A1(\mem[80] [2]), .A2(n_1_1_1138), .B1(n_1_1_1093), 
      .B2(\mem[34] [2]), .ZN(n_1_1_154));
   AOI221_X1 i_1_1_158 (.A(n_1_1_156), .B1(n_1_1_1072), .B2(\mem[6] [2]), 
      .C1(\mem[94] [2]), .C2(n_1_1_1157), .ZN(n_1_1_155));
   NAND3_X1 i_1_1_159 (.A1(n_1_1_190), .A2(n_1_1_168), .A3(n_1_1_157), .ZN(
      n_1_1_156));
   AOI22_X1 i_1_1_160 (.A1(\mem[93] [2]), .A2(n_1_1_1155), .B1(n_1_1_1041), 
      .B2(\mem[7] [2]), .ZN(n_1_1_157));
   NAND4_X1 i_1_1_161 (.A1(n_1_1_171), .A2(n_1_1_167), .A3(n_1_1_160), .A4(
      n_1_1_159), .ZN(n_1_1_158));
   AOI222_X1 i_1_1_162 (.A1(\mem[64] [2]), .A2(n_1_1_1118), .B1(n_1_1_1083), 
      .B2(\mem[24] [2]), .C1(n_1_1_1053), .C2(\mem[95] [2]), .ZN(n_1_1_159));
   AOI222_X1 i_1_1_163 (.A1(\mem[35] [2]), .A2(n_1_1_1094), .B1(n_1_1_1092), 
      .B2(\mem[33] [2]), .C1(n_1_1_1062), .C2(\mem[84] [2]), .ZN(n_1_1_160));
   AOI221_X1 i_1_1_164 (.A(n_1_1_162), .B1(n_1_1_1074), .B2(\mem[9] [2]), 
      .C1(\mem[21] [2]), .C2(n_1_1_1081), .ZN(n_1_1_161));
   NAND3_X1 i_1_1_165 (.A1(n_1_1_189), .A2(n_1_1_188), .A3(n_1_1_186), .ZN(
      n_1_1_162));
   AOI22_X1 i_1_1_166 (.A1(\mem[67] [2]), .A2(n_1_1_1121), .B1(n_1_1_1026), 
      .B2(\mem[56] [2]), .ZN(n_1_1_163));
   AOI222_X1 i_1_1_167 (.A1(\mem[3] [2]), .A2(n_1_1_1069), .B1(n_1_1_1063), 
      .B2(\mem[11] [2]), .C1(\mem[88] [2]), .C2(n_1_1_1056), .ZN(n_1_1_164));
   AOI22_X1 i_1_1_168 (.A1(\mem[87] [2]), .A2(n_1_1_1144), .B1(n_1_1_1134), 
      .B2(\mem[78] [2]), .ZN(n_1_1_165));
   AOI22_X1 i_1_1_169 (.A1(\mem[71] [2]), .A2(n_1_1_1126), .B1(n_1_1_1043), 
      .B2(\mem[53] [2]), .ZN(n_1_1_166));
   AOI22_X1 i_1_1_170 (.A1(\mem[26] [2]), .A2(n_1_1_1044), .B1(n_1_1_1040), 
      .B2(\mem[52] [2]), .ZN(n_1_1_167));
   AOI22_X1 i_1_1_171 (.A1(\mem[19] [2]), .A2(n_1_1_1080), .B1(n_1_1_1025), 
      .B2(\mem[43] [2]), .ZN(n_1_1_168));
   AOI22_X1 i_1_1_172 (.A1(\mem[81] [2]), .A2(n_1_1_1139), .B1(n_1_1_1123), 
      .B2(\mem[69] [2]), .ZN(n_1_1_169));
   AOI22_X1 i_1_1_173 (.A1(\mem[92] [2]), .A2(n_1_1_1153), .B1(n_1_1_1028), 
      .B2(\mem[82] [2]), .ZN(n_1_1_170));
   AOI221_X1 i_1_1_174 (.A(n_1_1_172), .B1(n_1_1_1097), .B2(\mem[38] [2]), 
      .C1(\mem[42] [2]), .C2(n_1_1_1033), .ZN(n_1_1_171));
   NAND3_X1 i_1_1_175 (.A1(n_1_1_182), .A2(n_1_1_174), .A3(n_1_1_173), .ZN(
      n_1_1_172));
   AOI22_X1 i_1_1_176 (.A1(\mem[25] [2]), .A2(n_1_1_1084), .B1(n_1_1_1078), 
      .B2(\mem[16] [2]), .ZN(n_1_1_173));
   AOI22_X1 i_1_1_177 (.A1(\mem[96] [2]), .A2(n_1_1_1163), .B1(n_1_1_1109), 
      .B2(\mem[58] [2]), .ZN(n_1_1_174));
   AOI22_X1 i_1_1_178 (.A1(\mem[55] [2]), .A2(n_1_1_1107), .B1(n_1_1_1031), 
      .B2(\mem[39] [2]), .ZN(n_1_1_175));
   AOI22_X1 i_1_1_179 (.A1(\mem[4] [2]), .A2(n_1_1_1070), .B1(n_1_1_1046), 
      .B2(\mem[60] [2]), .ZN(n_1_1_176));
   AOI22_X1 i_1_1_180 (.A1(\mem[41] [2]), .A2(n_1_1_1100), .B1(n_1_1_1096), 
      .B2(\mem[37] [2]), .ZN(n_1_1_177));
   AOI22_X1 i_1_1_181 (.A1(\mem[49] [2]), .A2(n_1_1_1105), .B1(n_1_1_1035), 
      .B2(\mem[50] [2]), .ZN(n_1_1_178));
   AOI22_X1 i_1_1_182 (.A1(\mem[8] [2]), .A2(n_1_1_1073), .B1(n_1_1_1039), 
      .B2(\mem[76] [2]), .ZN(n_1_1_179));
   AOI22_X1 i_1_1_183 (.A1(\mem[79] [2]), .A2(n_1_1_1135), .B1(n_1_1_1104), 
      .B2(\mem[48] [2]), .ZN(n_1_1_180));
   AOI22_X1 i_1_1_184 (.A1(\mem[1] [2]), .A2(n_1_1_1067), .B1(n_1_1_1029), 
      .B2(\mem[62] [2]), .ZN(n_1_1_181));
   AOI22_X1 i_1_1_185 (.A1(\mem[100] [2]), .A2(n_1_1_1174), .B1(n_1_1_1038), 
      .B2(\mem[15] [2]), .ZN(n_1_1_182));
   AOI22_X1 i_1_1_186 (.A1(\mem[97] [2]), .A2(n_1_1_1165), .B1(n_1_1_1036), 
      .B2(\mem[14] [2]), .ZN(n_1_1_183));
   AOI22_X1 i_1_1_187 (.A1(\mem[99] [2]), .A2(n_1_1_1171), .B1(n_1_1_1088), 
      .B2(\mem[31] [2]), .ZN(n_1_1_184));
   AOI22_X1 i_1_1_188 (.A1(\mem[98] [2]), .A2(n_1_1_1168), .B1(n_1_1_1068), 
      .B2(\mem[2] [2]), .ZN(n_1_1_185));
   AOI22_X1 i_1_1_189 (.A1(\mem[22] [2]), .A2(n_1_1_1054), .B1(n_1_1_1051), 
      .B2(\mem[29] [2]), .ZN(n_1_1_186));
   AOI22_X1 i_1_1_190 (.A1(\mem[77] [2]), .A2(n_1_1_1133), .B1(n_1_1_1071), 
      .B2(\mem[5] [2]), .ZN(n_1_1_187));
   AOI22_X1 i_1_1_191 (.A1(\mem[75] [2]), .A2(n_1_1_1061), .B1(n_1_1_1047), 
      .B2(\mem[83] [2]), .ZN(n_1_1_188));
   AOI22_X1 i_1_1_192 (.A1(\mem[54] [2]), .A2(n_1_1_1106), .B1(n_1_1_1030), 
      .B2(\mem[20] [2]), .ZN(n_1_1_189));
   AOI22_X1 i_1_1_193 (.A1(\mem[70] [2]), .A2(n_1_1_1125), .B1(n_1_1_1027), 
      .B2(\mem[27] [2]), .ZN(n_1_1_190));
   AOI22_X1 i_1_1_194 (.A1(\mem[40] [2]), .A2(n_1_1_1099), .B1(n_1_1_1058), 
      .B2(\mem[85] [2]), .ZN(n_1_1_191));
   NOR2_X1 i_1_1_195 (.A1(read_signal), .A2(dataout[2]), .ZN(n_1_1_192));
   MUX2_X1 i_1_1_196 (.A(dataout[3]), .B(n_1_1_193), .S(read_signal), .Z(n_1_3));
   NAND3_X1 i_1_1_197 (.A1(n_1_1_238), .A2(n_1_1_237), .A3(n_1_1_194), .ZN(
      n_1_1_193));
   NOR4_X1 i_1_1_198 (.A1(n_1_1_232), .A2(n_1_1_220), .A3(n_1_1_202), .A4(
      n_1_1_195), .ZN(n_1_1_194));
   NAND3_X1 i_1_1_199 (.A1(n_1_1_245), .A2(n_1_1_199), .A3(n_1_1_196), .ZN(
      n_1_1_195));
   AOI221_X1 i_1_1_200 (.A(n_1_1_197), .B1(n_1_1_1080), .B2(\mem[19] [3]), 
      .C1(\mem[33] [3]), .C2(n_1_1_1092), .ZN(n_1_1_196));
   NAND3_X1 i_1_1_201 (.A1(n_1_1_246), .A2(n_1_1_244), .A3(n_1_1_198), .ZN(
      n_1_1_197));
   AOI22_X1 i_1_1_202 (.A1(\mem[83] [3]), .A2(n_1_1_1047), .B1(n_1_1_1041), 
      .B2(\mem[7] [3]), .ZN(n_1_1_198));
   AOI221_X1 i_1_1_203 (.A(n_1_1_200), .B1(n_1_1_1042), .B2(\mem[12] [3]), 
      .C1(\mem[80] [3]), .C2(n_1_1_1138), .ZN(n_1_1_199));
   NAND3_X1 i_1_1_204 (.A1(n_1_1_248), .A2(n_1_1_247), .A3(n_1_1_201), .ZN(
      n_1_1_200));
   AOI22_X1 i_1_1_205 (.A1(\mem[63] [3]), .A2(n_1_1_1116), .B1(n_1_1_1083), 
      .B2(\mem[24] [3]), .ZN(n_1_1_201));
   NAND4_X1 i_1_1_206 (.A1(n_1_1_252), .A2(n_1_1_213), .A3(n_1_1_208), .A4(
      n_1_1_203), .ZN(n_1_1_202));
   AOI221_X1 i_1_1_207 (.A(n_1_1_204), .B1(n_1_1_1025), .B2(\mem[43] [3]), 
      .C1(\mem[98] [3]), .C2(n_1_1_1168), .ZN(n_1_1_203));
   NAND3_X1 i_1_1_208 (.A1(n_1_1_207), .A2(n_1_1_206), .A3(n_1_1_205), .ZN(
      n_1_1_204));
   AOI22_X1 i_1_1_209 (.A1(\mem[89] [3]), .A2(n_1_1_1148), .B1(n_1_1_1087), 
      .B2(\mem[30] [3]), .ZN(n_1_1_205));
   AOI222_X1 i_1_1_210 (.A1(\mem[13] [3]), .A2(n_1_1_1075), .B1(n_1_1_1069), 
      .B2(\mem[3] [3]), .C1(n_1_1_1046), .C2(\mem[60] [3]), .ZN(n_1_1_206));
   AOI22_X1 i_1_1_211 (.A1(\mem[74] [3]), .A2(n_1_1_1055), .B1(n_1_1_1039), 
      .B2(\mem[76] [3]), .ZN(n_1_1_207));
   AOI221_X1 i_1_1_212 (.A(n_1_1_209), .B1(n_1_1_1094), .B2(\mem[35] [3]), 
      .C1(\mem[52] [3]), .C2(n_1_1_1040), .ZN(n_1_1_208));
   NAND3_X1 i_1_1_213 (.A1(n_1_1_212), .A2(n_1_1_211), .A3(n_1_1_210), .ZN(
      n_1_1_209));
   AOI22_X1 i_1_1_214 (.A1(\mem[69] [3]), .A2(n_1_1_1123), .B1(n_1_1_1108), 
      .B2(\mem[57] [3]), .ZN(n_1_1_210));
   AOI22_X1 i_1_1_215 (.A1(\mem[79] [3]), .A2(n_1_1_1135), .B1(n_1_1_1105), 
      .B2(\mem[49] [3]), .ZN(n_1_1_211));
   AOI22_X1 i_1_1_216 (.A1(\mem[46] [3]), .A2(n_1_1_1101), .B1(n_1_1_1056), 
      .B2(\mem[88] [3]), .ZN(n_1_1_212));
   AOI211_X1 i_1_1_217 (.A(n_1_1_217), .B(n_1_1_214), .C1(\mem[9] [3]), .C2(
      n_1_1_1074), .ZN(n_1_1_213));
   NAND3_X1 i_1_1_218 (.A1(n_1_1_243), .A2(n_1_1_216), .A3(n_1_1_215), .ZN(
      n_1_1_214));
   AOI222_X1 i_1_1_219 (.A1(\mem[99] [3]), .A2(n_1_1_1171), .B1(n_1_1_1097), 
      .B2(\mem[38] [3]), .C1(n_1_1_1088), .C2(\mem[31] [3]), .ZN(n_1_1_215));
   AOI22_X1 i_1_1_220 (.A1(\mem[64] [3]), .A2(n_1_1_1118), .B1(n_1_1_1111), 
      .B2(\mem[59] [3]), .ZN(n_1_1_216));
   NAND4_X1 i_1_1_221 (.A1(n_1_1_253), .A2(n_1_1_218), .A3(n_1_1_249), .A4(
      n_1_1_219), .ZN(n_1_1_217));
   AOI222_X1 i_1_1_222 (.A1(\mem[73] [3]), .A2(n_1_1_1129), .B1(n_1_1_1070), 
      .B2(\mem[4] [3]), .C1(n_1_1_1029), .C2(\mem[62] [3]), .ZN(n_1_1_218));
   AOI22_X1 i_1_1_223 (.A1(\mem[68] [3]), .A2(n_1_1_1122), .B1(n_1_1_1064), 
      .B2(\mem[18] [3]), .ZN(n_1_1_219));
   NAND4_X1 i_1_1_224 (.A1(n_1_1_231), .A2(n_1_1_230), .A3(n_1_1_226), .A4(
      n_1_1_221), .ZN(n_1_1_220));
   AOI221_X1 i_1_1_225 (.A(n_1_1_222), .B1(n_1_1_1067), .B2(\mem[1] [3]), 
      .C1(\mem[5] [3]), .C2(n_1_1_1071), .ZN(n_1_1_221));
   NAND4_X1 i_1_1_226 (.A1(n_1_1_250), .A2(n_1_1_225), .A3(n_1_1_224), .A4(
      n_1_1_223), .ZN(n_1_1_222));
   AOI22_X1 i_1_1_227 (.A1(\mem[41] [3]), .A2(n_1_1_1100), .B1(n_1_1_1048), 
      .B2(\mem[10] [3]), .ZN(n_1_1_223));
   AOI22_X1 i_1_1_228 (.A1(\mem[67] [3]), .A2(n_1_1_1121), .B1(n_1_1_1060), 
      .B2(\mem[28] [3]), .ZN(n_1_1_224));
   AOI22_X1 i_1_1_229 (.A1(\mem[77] [3]), .A2(n_1_1_1133), .B1(n_1_1_1072), 
      .B2(\mem[6] [3]), .ZN(n_1_1_225));
   AOI221_X1 i_1_1_230 (.A(n_1_1_227), .B1(n_1_1_1061), .B2(\mem[75] [3]), 
      .C1(\mem[90] [3]), .C2(n_1_1_1050), .ZN(n_1_1_226));
   NAND3_X1 i_1_1_231 (.A1(n_1_1_251), .A2(n_1_1_229), .A3(n_1_1_228), .ZN(
      n_1_1_227));
   AOI22_X1 i_1_1_232 (.A1(\mem[53] [3]), .A2(n_1_1_1043), .B1(n_1_1_1026), 
      .B2(\mem[56] [3]), .ZN(n_1_1_228));
   AOI22_X1 i_1_1_233 (.A1(\mem[96] [3]), .A2(n_1_1_1163), .B1(n_1_1_1044), 
      .B2(\mem[26] [3]), .ZN(n_1_1_229));
   AOI222_X1 i_1_1_234 (.A1(\mem[100] [3]), .A2(n_1_1_1174), .B1(n_1_1_1165), 
      .B2(\mem[97] [3]), .C1(n_1_1_1054), .C2(\mem[22] [3]), .ZN(n_1_1_230));
   AOI222_X1 i_1_1_235 (.A1(\mem[85] [3]), .A2(n_1_1_1058), .B1(n_1_1_1057), 
      .B2(\mem[61] [3]), .C1(\mem[11] [3]), .C2(n_1_1_1063), .ZN(n_1_1_231));
   NAND4_X1 i_1_1_236 (.A1(n_1_1_236), .A2(n_1_1_235), .A3(n_1_1_234), .A4(
      n_1_1_233), .ZN(n_1_1_232));
   AOI22_X1 i_1_1_237 (.A1(\mem[93] [3]), .A2(n_1_1_1155), .B1(n_1_1_1059), 
      .B2(\mem[51] [3]), .ZN(n_1_1_233));
   AOI22_X1 i_1_1_238 (.A1(\mem[2] [3]), .A2(n_1_1_1068), .B1(n_1_1_1051), 
      .B2(\mem[29] [3]), .ZN(n_1_1_234));
   AOI222_X1 i_1_1_239 (.A1(\mem[54] [3]), .A2(n_1_1_1106), .B1(n_1_1_1104), 
      .B2(\mem[48] [3]), .C1(n_1_1_1030), .C2(\mem[20] [3]), .ZN(n_1_1_235));
   AOI222_X1 i_1_1_240 (.A1(\mem[94] [3]), .A2(n_1_1_1157), .B1(n_1_1_1081), 
      .B2(\mem[21] [3]), .C1(n_1_1_1032), .C2(\mem[44] [3]), .ZN(n_1_1_236));
   AOI222_X1 i_1_1_241 (.A1(\mem[87] [3]), .A2(n_1_1_1144), .B1(n_1_1_1134), 
      .B2(\mem[78] [3]), .C1(n_1_1_1062), .C2(\mem[84] [3]), .ZN(n_1_1_237));
   AOI221_X1 i_1_1_242 (.A(n_1_1_239), .B1(n_1_1_1078), .B2(\mem[16] [3]), 
      .C1(\mem[42] [3]), .C2(n_1_1_1033), .ZN(n_1_1_238));
   NAND3_X1 i_1_1_243 (.A1(n_1_1_242), .A2(n_1_1_241), .A3(n_1_1_240), .ZN(
      n_1_1_239));
   AOI222_X1 i_1_1_244 (.A1(\mem[65] [3]), .A2(n_1_1_1119), .B1(n_1_1_1109), 
      .B2(\mem[58] [3]), .C1(n_1_1_1037), .C2(\mem[91] [3]), .ZN(n_1_1_240));
   AOI222_X1 i_1_1_245 (.A1(\mem[70] [3]), .A2(n_1_1_1125), .B1(n_1_1_1084), 
      .B2(\mem[25] [3]), .C1(n_1_1_1045), .C2(\mem[45] [3]), .ZN(n_1_1_241));
   AOI222_X1 i_1_1_246 (.A1(\mem[86] [3]), .A2(n_1_1_1142), .B1(n_1_1_1099), 
      .B2(\mem[40] [3]), .C1(n_1_1_1038), .C2(\mem[15] [3]), .ZN(n_1_1_242));
   AOI22_X1 i_1_1_247 (.A1(\mem[66] [3]), .A2(n_1_1_1120), .B1(n_1_1_1036), 
      .B2(\mem[14] [3]), .ZN(n_1_1_243));
   AOI22_X1 i_1_1_248 (.A1(\mem[72] [3]), .A2(n_1_1_1127), .B1(n_1_1_1027), 
      .B2(\mem[27] [3]), .ZN(n_1_1_244));
   AOI22_X1 i_1_1_249 (.A1(\mem[95] [3]), .A2(n_1_1_1053), .B1(n_1_1_1052), 
      .B2(\mem[23] [3]), .ZN(n_1_1_245));
   AOI22_X1 i_1_1_250 (.A1(\mem[81] [3]), .A2(n_1_1_1139), .B1(n_1_1_1066), 
      .B2(\mem[0] [3]), .ZN(n_1_1_246));
   AOI22_X1 i_1_1_251 (.A1(\mem[36] [3]), .A2(n_1_1_1095), .B1(n_1_1_1049), 
      .B2(\mem[17] [3]), .ZN(n_1_1_247));
   AOI22_X1 i_1_1_252 (.A1(\mem[71] [3]), .A2(n_1_1_1126), .B1(n_1_1_1102), 
      .B2(\mem[47] [3]), .ZN(n_1_1_248));
   NAND2_X1 i_1_1_253 (.A1(\mem[37] [3]), .A2(n_1_1_1096), .ZN(n_1_1_249));
   AOI22_X1 i_1_1_254 (.A1(\mem[34] [3]), .A2(n_1_1_1093), .B1(n_1_1_1073), 
      .B2(\mem[8] [3]), .ZN(n_1_1_250));
   AOI22_X1 i_1_1_255 (.A1(\mem[92] [3]), .A2(n_1_1_1153), .B1(n_1_1_1028), 
      .B2(\mem[82] [3]), .ZN(n_1_1_251));
   AOI22_X1 i_1_1_256 (.A1(\mem[32] [3]), .A2(n_1_1_1091), .B1(n_1_1_1035), 
      .B2(\mem[50] [3]), .ZN(n_1_1_252));
   AOI22_X1 i_1_1_257 (.A1(\mem[55] [3]), .A2(n_1_1_1107), .B1(n_1_1_1031), 
      .B2(\mem[39] [3]), .ZN(n_1_1_253));
   AOI21_X1 i_1_1_258 (.A(n_1_1_254), .B1(n_1_1_255), .B2(n_1_1_287), .ZN(n_1_4));
   NOR2_X1 i_1_1_259 (.A1(read_signal), .A2(dataout[4]), .ZN(n_1_1_254));
   NOR4_X1 i_1_1_260 (.A1(n_1_1_282), .A2(n_1_1_278), .A3(n_1_1_258), .A4(
      n_1_1_256), .ZN(n_1_1_255));
   NAND4_X1 i_1_1_261 (.A1(read_signal), .A2(n_1_1_318), .A3(n_1_1_315), 
      .A4(n_1_1_257), .ZN(n_1_1_256));
   AOI22_X1 i_1_1_262 (.A1(\mem[37] [4]), .A2(n_1_1_1096), .B1(n_1_1_1057), 
      .B2(\mem[61] [4]), .ZN(n_1_1_257));
   NAND4_X1 i_1_1_263 (.A1(n_1_1_273), .A2(n_1_1_268), .A3(n_1_1_263), .A4(
      n_1_1_259), .ZN(n_1_1_258));
   AOI221_X1 i_1_1_264 (.A(n_1_1_260), .B1(n_1_1_1081), .B2(\mem[21] [4]), 
      .C1(\mem[80] [4]), .C2(n_1_1_1138), .ZN(n_1_1_259));
   NAND3_X1 i_1_1_265 (.A1(n_1_1_316), .A2(n_1_1_262), .A3(n_1_1_261), .ZN(
      n_1_1_260));
   AOI22_X1 i_1_1_266 (.A1(\mem[70] [4]), .A2(n_1_1_1125), .B1(n_1_1_1033), 
      .B2(\mem[42] [4]), .ZN(n_1_1_261));
   AOI22_X1 i_1_1_267 (.A1(\mem[30] [4]), .A2(n_1_1_1087), .B1(n_1_1_1044), 
      .B2(\mem[26] [4]), .ZN(n_1_1_262));
   AOI221_X1 i_1_1_268 (.A(n_1_1_264), .B1(n_1_1_1097), .B2(\mem[38] [4]), 
      .C1(\mem[48] [4]), .C2(n_1_1_1104), .ZN(n_1_1_263));
   NAND3_X1 i_1_1_269 (.A1(n_1_1_267), .A2(n_1_1_266), .A3(n_1_1_265), .ZN(
      n_1_1_264));
   AOI22_X1 i_1_1_270 (.A1(\mem[100] [4]), .A2(n_1_1_1174), .B1(n_1_1_1029), 
      .B2(\mem[62] [4]), .ZN(n_1_1_265));
   AOI22_X1 i_1_1_271 (.A1(\mem[2] [4]), .A2(n_1_1_1068), .B1(n_1_1_1041), 
      .B2(\mem[7] [4]), .ZN(n_1_1_266));
   AOI22_X1 i_1_1_272 (.A1(\mem[94] [4]), .A2(n_1_1_1157), .B1(n_1_1_1025), 
      .B2(\mem[43] [4]), .ZN(n_1_1_267));
   AOI221_X1 i_1_1_273 (.A(n_1_1_269), .B1(n_1_1_1102), .B2(\mem[47] [4]), 
      .C1(\mem[75] [4]), .C2(n_1_1_1061), .ZN(n_1_1_268));
   NAND3_X1 i_1_1_274 (.A1(n_1_1_272), .A2(n_1_1_271), .A3(n_1_1_270), .ZN(
      n_1_1_269));
   AOI22_X1 i_1_1_275 (.A1(\mem[28] [4]), .A2(n_1_1_1060), .B1(n_1_1_1035), 
      .B2(\mem[50] [4]), .ZN(n_1_1_270));
   AOI22_X1 i_1_1_276 (.A1(\mem[33] [4]), .A2(n_1_1_1092), .B1(n_1_1_1053), 
      .B2(\mem[95] [4]), .ZN(n_1_1_271));
   AOI22_X1 i_1_1_277 (.A1(\mem[54] [4]), .A2(n_1_1_1106), .B1(n_1_1_1030), 
      .B2(\mem[20] [4]), .ZN(n_1_1_272));
   AOI221_X1 i_1_1_278 (.A(n_1_1_274), .B1(n_1_1_1049), .B2(\mem[17] [4]), 
      .C1(\mem[96] [4]), .C2(n_1_1_1163), .ZN(n_1_1_273));
   NAND3_X1 i_1_1_279 (.A1(n_1_1_277), .A2(n_1_1_276), .A3(n_1_1_275), .ZN(
      n_1_1_274));
   AOI22_X1 i_1_1_280 (.A1(\mem[65] [4]), .A2(n_1_1_1119), .B1(n_1_1_1032), 
      .B2(\mem[44] [4]), .ZN(n_1_1_275));
   AOI22_X1 i_1_1_281 (.A1(\mem[97] [4]), .A2(n_1_1_1165), .B1(n_1_1_1071), 
      .B2(\mem[5] [4]), .ZN(n_1_1_276));
   AOI22_X1 i_1_1_282 (.A1(\mem[72] [4]), .A2(n_1_1_1127), .B1(n_1_1_1093), 
      .B2(\mem[34] [4]), .ZN(n_1_1_277));
   NAND4_X1 i_1_1_283 (.A1(n_1_1_317), .A2(n_1_1_281), .A3(n_1_1_280), .A4(
      n_1_1_279), .ZN(n_1_1_278));
   AOI22_X1 i_1_1_284 (.A1(\mem[51] [4]), .A2(n_1_1_1059), .B1(n_1_1_1054), 
      .B2(\mem[22] [4]), .ZN(n_1_1_279));
   AOI22_X1 i_1_1_285 (.A1(\mem[63] [4]), .A2(n_1_1_1116), .B1(n_1_1_1101), 
      .B2(\mem[46] [4]), .ZN(n_1_1_280));
   AOI22_X1 i_1_1_286 (.A1(\mem[6] [4]), .A2(n_1_1_1072), .B1(n_1_1_1036), 
      .B2(\mem[14] [4]), .ZN(n_1_1_281));
   NAND4_X1 i_1_1_287 (.A1(n_1_1_286), .A2(n_1_1_285), .A3(n_1_1_284), .A4(
      n_1_1_283), .ZN(n_1_1_282));
   AOI22_X1 i_1_1_288 (.A1(\mem[1] [4]), .A2(n_1_1_1067), .B1(n_1_1_1038), 
      .B2(\mem[15] [4]), .ZN(n_1_1_283));
   AOI22_X1 i_1_1_289 (.A1(\mem[19] [4]), .A2(n_1_1_1080), .B1(n_1_1_1063), 
      .B2(\mem[11] [4]), .ZN(n_1_1_284));
   AOI22_X1 i_1_1_290 (.A1(\mem[18] [4]), .A2(n_1_1_1064), .B1(n_1_1_1027), 
      .B2(\mem[27] [4]), .ZN(n_1_1_285));
   AOI22_X1 i_1_1_291 (.A1(\mem[92] [4]), .A2(n_1_1_1153), .B1(n_1_1_1083), 
      .B2(\mem[24] [4]), .ZN(n_1_1_286));
   NOR3_X1 i_1_1_292 (.A1(n_1_1_309), .A2(n_1_1_302), .A3(n_1_1_288), .ZN(
      n_1_1_287));
   NAND3_X1 i_1_1_293 (.A1(n_1_1_297), .A2(n_1_1_293), .A3(n_1_1_289), .ZN(
      n_1_1_288));
   AOI221_X1 i_1_1_294 (.A(n_1_1_290), .B1(n_1_1_1070), .B2(\mem[4] [4]), 
      .C1(\mem[52] [4]), .C2(n_1_1_1040), .ZN(n_1_1_289));
   NAND3_X1 i_1_1_295 (.A1(n_1_1_319), .A2(n_1_1_292), .A3(n_1_1_291), .ZN(
      n_1_1_290));
   AOI22_X1 i_1_1_296 (.A1(\mem[68] [4]), .A2(n_1_1_1122), .B1(n_1_1_1043), 
      .B2(\mem[53] [4]), .ZN(n_1_1_291));
   AOI22_X1 i_1_1_297 (.A1(\mem[86] [4]), .A2(n_1_1_1142), .B1(n_1_1_1075), 
      .B2(\mem[13] [4]), .ZN(n_1_1_292));
   AOI221_X1 i_1_1_298 (.A(n_1_1_294), .B1(n_1_1_1074), .B2(\mem[9] [4]), 
      .C1(\mem[98] [4]), .C2(n_1_1_1168), .ZN(n_1_1_293));
   NAND3_X1 i_1_1_299 (.A1(n_1_1_320), .A2(n_1_1_296), .A3(n_1_1_295), .ZN(
      n_1_1_294));
   AOI22_X1 i_1_1_300 (.A1(\mem[71] [4]), .A2(n_1_1_1126), .B1(n_1_1_1050), 
      .B2(\mem[90] [4]), .ZN(n_1_1_295));
   AOI22_X1 i_1_1_301 (.A1(\mem[57] [4]), .A2(n_1_1_1108), .B1(n_1_1_1095), 
      .B2(\mem[36] [4]), .ZN(n_1_1_296));
   AOI221_X1 i_1_1_302 (.A(n_1_1_298), .B1(n_1_1_1052), .B2(\mem[23] [4]), 
      .C1(\mem[87] [4]), .C2(n_1_1_1144), .ZN(n_1_1_297));
   NAND3_X1 i_1_1_303 (.A1(n_1_1_301), .A2(n_1_1_300), .A3(n_1_1_299), .ZN(
      n_1_1_298));
   AOI22_X1 i_1_1_304 (.A1(\mem[78] [4]), .A2(n_1_1_1134), .B1(n_1_1_1133), 
      .B2(\mem[77] [4]), .ZN(n_1_1_299));
   AOI22_X1 i_1_1_305 (.A1(\mem[85] [4]), .A2(n_1_1_1058), .B1(n_1_1_1039), 
      .B2(\mem[76] [4]), .ZN(n_1_1_300));
   AOI22_X1 i_1_1_306 (.A1(\mem[79] [4]), .A2(n_1_1_1135), .B1(n_1_1_1055), 
      .B2(\mem[74] [4]), .ZN(n_1_1_301));
   NAND4_X1 i_1_1_307 (.A1(n_1_1_321), .A2(n_1_1_314), .A3(n_1_1_304), .A4(
      n_1_1_303), .ZN(n_1_1_302));
   AOI222_X1 i_1_1_308 (.A1(\mem[89] [4]), .A2(n_1_1_1148), .B1(n_1_1_1111), 
      .B2(\mem[59] [4]), .C1(n_1_1_1073), .C2(\mem[8] [4]), .ZN(n_1_1_303));
   AOI221_X1 i_1_1_309 (.A(n_1_1_305), .B1(n_1_1_1139), .B2(\mem[81] [4]), 
      .C1(\mem[82] [4]), .C2(n_1_1_1028), .ZN(n_1_1_304));
   NAND3_X1 i_1_1_310 (.A1(n_1_1_308), .A2(n_1_1_307), .A3(n_1_1_306), .ZN(
      n_1_1_305));
   AOI22_X1 i_1_1_311 (.A1(\mem[73] [4]), .A2(n_1_1_1129), .B1(n_1_1_1051), 
      .B2(\mem[29] [4]), .ZN(n_1_1_306));
   AOI22_X1 i_1_1_312 (.A1(\mem[25] [4]), .A2(n_1_1_1084), .B1(n_1_1_1045), 
      .B2(\mem[45] [4]), .ZN(n_1_1_307));
   AOI22_X1 i_1_1_313 (.A1(\mem[12] [4]), .A2(n_1_1_1042), .B1(n_1_1_1037), 
      .B2(\mem[91] [4]), .ZN(n_1_1_308));
   NAND4_X1 i_1_1_314 (.A1(n_1_1_313), .A2(n_1_1_312), .A3(n_1_1_311), .A4(
      n_1_1_310), .ZN(n_1_1_309));
   AOI22_X1 i_1_1_315 (.A1(\mem[3] [4]), .A2(n_1_1_1069), .B1(n_1_1_1062), 
      .B2(\mem[84] [4]), .ZN(n_1_1_310));
   AOI22_X1 i_1_1_316 (.A1(\mem[69] [4]), .A2(n_1_1_1123), .B1(n_1_1_1088), 
      .B2(\mem[31] [4]), .ZN(n_1_1_311));
   AOI22_X1 i_1_1_317 (.A1(\mem[99] [4]), .A2(n_1_1_1171), .B1(n_1_1_1066), 
      .B2(\mem[0] [4]), .ZN(n_1_1_312));
   AOI22_X1 i_1_1_318 (.A1(\mem[93] [4]), .A2(n_1_1_1155), .B1(n_1_1_1105), 
      .B2(\mem[49] [4]), .ZN(n_1_1_313));
   AOI222_X1 i_1_1_319 (.A1(\mem[67] [4]), .A2(n_1_1_1121), .B1(n_1_1_1048), 
      .B2(\mem[10] [4]), .C1(n_1_1_1056), .C2(\mem[88] [4]), .ZN(n_1_1_314));
   NAND2_X1 i_1_1_320 (.A1(\mem[16] [4]), .A2(n_1_1_1078), .ZN(n_1_1_315));
   AOI22_X1 i_1_1_321 (.A1(\mem[58] [4]), .A2(n_1_1_1109), .B1(n_1_1_1047), 
      .B2(\mem[83] [4]), .ZN(n_1_1_316));
   AOI22_X1 i_1_1_322 (.A1(\mem[66] [4]), .A2(n_1_1_1120), .B1(n_1_1_1100), 
      .B2(\mem[41] [4]), .ZN(n_1_1_317));
   AOI22_X1 i_1_1_323 (.A1(\mem[55] [4]), .A2(n_1_1_1107), .B1(n_1_1_1099), 
      .B2(\mem[40] [4]), .ZN(n_1_1_318));
   AOI22_X1 i_1_1_324 (.A1(\mem[39] [4]), .A2(n_1_1_1031), .B1(n_1_1_1026), 
      .B2(\mem[56] [4]), .ZN(n_1_1_319));
   AOI22_X1 i_1_1_325 (.A1(\mem[32] [4]), .A2(n_1_1_1091), .B1(n_1_1_1046), 
      .B2(\mem[60] [4]), .ZN(n_1_1_320));
   AOI22_X1 i_1_1_326 (.A1(\mem[64] [4]), .A2(n_1_1_1118), .B1(n_1_1_1094), 
      .B2(\mem[35] [4]), .ZN(n_1_1_321));
   MUX2_X1 i_1_1_327 (.A(dataout[5]), .B(n_1_1_322), .S(read_signal), .Z(n_1_5));
   NAND4_X1 i_1_1_328 (.A1(n_1_1_350), .A2(n_1_1_327), .A3(n_1_1_324), .A4(
      n_1_1_323), .ZN(n_1_1_322));
   AOI221_X1 i_1_1_329 (.A(n_1_1_371), .B1(n_1_1_1045), .B2(\mem[45] [5]), 
      .C1(\mem[47] [5]), .C2(n_1_1_1102), .ZN(n_1_1_323));
   AOI221_X1 i_1_1_330 (.A(n_1_1_325), .B1(n_1_1_1091), .B2(\mem[32] [5]), 
      .C1(\mem[74] [5]), .C2(n_1_1_1055), .ZN(n_1_1_324));
   NAND3_X1 i_1_1_331 (.A1(n_1_1_383), .A2(n_1_1_380), .A3(n_1_1_326), .ZN(
      n_1_1_325));
   AOI22_X1 i_1_1_332 (.A1(\mem[100] [5]), .A2(n_1_1_1174), .B1(n_1_1_1056), 
      .B2(\mem[88] [5]), .ZN(n_1_1_326));
   AND4_X1 i_1_1_333 (.A1(n_1_1_368), .A2(n_1_1_331), .A3(n_1_1_330), .A4(
      n_1_1_328), .ZN(n_1_1_327));
   AOI221_X1 i_1_1_334 (.A(n_1_1_329), .B1(n_1_1_1105), .B2(\mem[49] [5]), 
      .C1(\mem[99] [5]), .C2(n_1_1_1171), .ZN(n_1_1_328));
   NAND3_X1 i_1_1_335 (.A1(n_1_1_370), .A2(n_1_1_369), .A3(n_1_1_367), .ZN(
      n_1_1_329));
   AOI222_X1 i_1_1_336 (.A1(\mem[25] [5]), .A2(n_1_1_1084), .B1(n_1_1_1074), 
      .B2(\mem[9] [5]), .C1(n_1_1_1060), .C2(\mem[28] [5]), .ZN(n_1_1_330));
   NOR4_X1 i_1_1_337 (.A1(n_1_1_345), .A2(n_1_1_341), .A3(n_1_1_337), .A4(
      n_1_1_332), .ZN(n_1_1_331));
   NAND4_X1 i_1_1_338 (.A1(n_1_1_336), .A2(n_1_1_335), .A3(n_1_1_334), .A4(
      n_1_1_333), .ZN(n_1_1_332));
   AOI22_X1 i_1_1_339 (.A1(\mem[81] [5]), .A2(n_1_1_1139), .B1(n_1_1_1129), 
      .B2(\mem[73] [5]), .ZN(n_1_1_333));
   AOI22_X1 i_1_1_340 (.A1(\mem[55] [5]), .A2(n_1_1_1107), .B1(n_1_1_1066), 
      .B2(\mem[0] [5]), .ZN(n_1_1_334));
   AOI22_X1 i_1_1_341 (.A1(\mem[84] [5]), .A2(n_1_1_1062), .B1(n_1_1_1044), 
      .B2(\mem[26] [5]), .ZN(n_1_1_335));
   AOI22_X1 i_1_1_342 (.A1(\mem[96] [5]), .A2(n_1_1_1163), .B1(n_1_1_1039), 
      .B2(\mem[76] [5]), .ZN(n_1_1_336));
   NAND4_X1 i_1_1_343 (.A1(n_1_1_382), .A2(n_1_1_340), .A3(n_1_1_339), .A4(
      n_1_1_338), .ZN(n_1_1_337));
   AOI22_X1 i_1_1_344 (.A1(\mem[48] [5]), .A2(n_1_1_1104), .B1(n_1_1_1041), 
      .B2(\mem[7] [5]), .ZN(n_1_1_338));
   AOI22_X1 i_1_1_345 (.A1(\mem[86] [5]), .A2(n_1_1_1142), .B1(n_1_1_1073), 
      .B2(\mem[8] [5]), .ZN(n_1_1_339));
   AOI22_X1 i_1_1_346 (.A1(\mem[33] [5]), .A2(n_1_1_1092), .B1(n_1_1_1081), 
      .B2(\mem[21] [5]), .ZN(n_1_1_340));
   NAND4_X1 i_1_1_347 (.A1(n_1_1_381), .A2(n_1_1_344), .A3(n_1_1_343), .A4(
      n_1_1_342), .ZN(n_1_1_341));
   AOI22_X1 i_1_1_348 (.A1(\mem[87] [5]), .A2(n_1_1_1144), .B1(n_1_1_1038), 
      .B2(\mem[15] [5]), .ZN(n_1_1_342));
   AOI22_X1 i_1_1_349 (.A1(\mem[19] [5]), .A2(n_1_1_1080), .B1(n_1_1_1033), 
      .B2(\mem[42] [5]), .ZN(n_1_1_343));
   AOI22_X1 i_1_1_350 (.A1(\mem[67] [5]), .A2(n_1_1_1121), .B1(n_1_1_1075), 
      .B2(\mem[13] [5]), .ZN(n_1_1_344));
   NAND4_X1 i_1_1_351 (.A1(n_1_1_349), .A2(n_1_1_348), .A3(n_1_1_347), .A4(
      n_1_1_346), .ZN(n_1_1_345));
   AOI22_X1 i_1_1_352 (.A1(\mem[2] [5]), .A2(n_1_1_1068), .B1(n_1_1_1057), 
      .B2(\mem[61] [5]), .ZN(n_1_1_346));
   AOI22_X1 i_1_1_353 (.A1(\mem[66] [5]), .A2(n_1_1_1120), .B1(n_1_1_1051), 
      .B2(\mem[29] [5]), .ZN(n_1_1_347));
   AOI22_X1 i_1_1_354 (.A1(\mem[36] [5]), .A2(n_1_1_1095), .B1(n_1_1_1036), 
      .B2(\mem[14] [5]), .ZN(n_1_1_348));
   AOI22_X1 i_1_1_355 (.A1(\mem[54] [5]), .A2(n_1_1_1106), .B1(n_1_1_1029), 
      .B2(\mem[62] [5]), .ZN(n_1_1_349));
   AND4_X1 i_1_1_356 (.A1(n_1_1_358), .A2(n_1_1_353), .A3(n_1_1_352), .A4(
      n_1_1_351), .ZN(n_1_1_350));
   AOI222_X1 i_1_1_357 (.A1(\mem[53] [5]), .A2(n_1_1_1043), .B1(n_1_1_1040), 
      .B2(\mem[52] [5]), .C1(\mem[37] [5]), .C2(n_1_1_1096), .ZN(n_1_1_351));
   AOI222_X1 i_1_1_358 (.A1(\mem[78] [5]), .A2(n_1_1_1134), .B1(n_1_1_1118), 
      .B2(\mem[64] [5]), .C1(n_1_1_1101), .C2(\mem[46] [5]), .ZN(n_1_1_352));
   AOI221_X1 i_1_1_359 (.A(n_1_1_354), .B1(n_1_1_1052), .B2(\mem[23] [5]), 
      .C1(\mem[44] [5]), .C2(n_1_1_1032), .ZN(n_1_1_353));
   NAND3_X1 i_1_1_360 (.A1(n_1_1_357), .A2(n_1_1_356), .A3(n_1_1_355), .ZN(
      n_1_1_354));
   AOI22_X1 i_1_1_361 (.A1(\mem[4] [5]), .A2(n_1_1_1070), .B1(n_1_1_1058), 
      .B2(\mem[85] [5]), .ZN(n_1_1_355));
   AOI22_X1 i_1_1_362 (.A1(\mem[68] [5]), .A2(n_1_1_1122), .B1(n_1_1_1111), 
      .B2(\mem[59] [5]), .ZN(n_1_1_356));
   AOI22_X1 i_1_1_363 (.A1(\mem[31] [5]), .A2(n_1_1_1088), .B1(n_1_1_1047), 
      .B2(\mem[83] [5]), .ZN(n_1_1_357));
   AOI221_X1 i_1_1_364 (.A(n_1_1_359), .B1(n_1_1_1042), .B2(\mem[12] [5]), 
      .C1(\mem[35] [5]), .C2(n_1_1_1094), .ZN(n_1_1_358));
   NAND4_X1 i_1_1_365 (.A1(n_1_1_366), .A2(n_1_1_362), .A3(n_1_1_361), .A4(
      n_1_1_360), .ZN(n_1_1_359));
   AOI22_X1 i_1_1_366 (.A1(\mem[91] [5]), .A2(n_1_1_1037), .B1(n_1_1_1025), 
      .B2(\mem[43] [5]), .ZN(n_1_1_360));
   AOI22_X1 i_1_1_367 (.A1(\mem[94] [5]), .A2(n_1_1_1157), .B1(n_1_1_1087), 
      .B2(\mem[30] [5]), .ZN(n_1_1_361));
   AOI221_X1 i_1_1_368 (.A(n_1_1_363), .B1(n_1_1_1069), .B2(\mem[3] [5]), 
      .C1(\mem[79] [5]), .C2(n_1_1_1135), .ZN(n_1_1_362));
   NAND3_X1 i_1_1_369 (.A1(n_1_1_384), .A2(n_1_1_365), .A3(n_1_1_364), .ZN(
      n_1_1_363));
   AOI22_X1 i_1_1_370 (.A1(\mem[51] [5]), .A2(n_1_1_1059), .B1(n_1_1_1046), 
      .B2(\mem[60] [5]), .ZN(n_1_1_364));
   AOI22_X1 i_1_1_371 (.A1(\mem[39] [5]), .A2(n_1_1_1031), .B1(n_1_1_1030), 
      .B2(\mem[20] [5]), .ZN(n_1_1_365));
   AOI22_X1 i_1_1_372 (.A1(\mem[77] [5]), .A2(n_1_1_1133), .B1(n_1_1_1064), 
      .B2(\mem[18] [5]), .ZN(n_1_1_366));
   AOI22_X1 i_1_1_373 (.A1(\mem[65] [5]), .A2(n_1_1_1119), .B1(n_1_1_1063), 
      .B2(\mem[11] [5]), .ZN(n_1_1_367));
   AOI22_X1 i_1_1_374 (.A1(\mem[63] [5]), .A2(n_1_1_1116), .B1(n_1_1_1099), 
      .B2(\mem[40] [5]), .ZN(n_1_1_368));
   AOI22_X1 i_1_1_375 (.A1(\mem[80] [5]), .A2(n_1_1_1138), .B1(n_1_1_1123), 
      .B2(\mem[69] [5]), .ZN(n_1_1_369));
   AOI22_X1 i_1_1_376 (.A1(\mem[16] [5]), .A2(n_1_1_1078), .B1(n_1_1_1027), 
      .B2(\mem[27] [5]), .ZN(n_1_1_370));
   NAND4_X1 i_1_1_377 (.A1(n_1_1_378), .A2(n_1_1_377), .A3(n_1_1_376), .A4(
      n_1_1_372), .ZN(n_1_1_371));
   AOI221_X1 i_1_1_378 (.A(n_1_1_373), .B1(n_1_1_1049), .B2(\mem[17] [5]), 
      .C1(\mem[56] [5]), .C2(n_1_1_1026), .ZN(n_1_1_372));
   NAND3_X1 i_1_1_379 (.A1(n_1_1_379), .A2(n_1_1_375), .A3(n_1_1_374), .ZN(
      n_1_1_373));
   AOI22_X1 i_1_1_380 (.A1(\mem[58] [5]), .A2(n_1_1_1109), .B1(n_1_1_1071), 
      .B2(\mem[5] [5]), .ZN(n_1_1_374));
   AOI22_X1 i_1_1_381 (.A1(\mem[34] [5]), .A2(n_1_1_1093), .B1(n_1_1_1048), 
      .B2(\mem[10] [5]), .ZN(n_1_1_375));
   AOI22_X1 i_1_1_382 (.A1(\mem[95] [5]), .A2(n_1_1_1053), .B1(n_1_1_1050), 
      .B2(\mem[90] [5]), .ZN(n_1_1_376));
   AOI222_X1 i_1_1_383 (.A1(\mem[71] [5]), .A2(n_1_1_1126), .B1(n_1_1_1035), 
      .B2(\mem[50] [5]), .C1(n_1_1_1028), .C2(\mem[82] [5]), .ZN(n_1_1_377));
   AOI222_X1 i_1_1_384 (.A1(\mem[38] [5]), .A2(n_1_1_1097), .B1(n_1_1_1054), 
      .B2(\mem[22] [5]), .C1(n_1_1_1061), .C2(\mem[75] [5]), .ZN(n_1_1_378));
   AOI22_X1 i_1_1_385 (.A1(\mem[97] [5]), .A2(n_1_1_1165), .B1(n_1_1_1083), 
      .B2(\mem[24] [5]), .ZN(n_1_1_379));
   AOI22_X1 i_1_1_386 (.A1(\mem[89] [5]), .A2(n_1_1_1148), .B1(n_1_1_1072), 
      .B2(\mem[6] [5]), .ZN(n_1_1_380));
   AOI22_X1 i_1_1_387 (.A1(\mem[41] [5]), .A2(n_1_1_1100), .B1(n_1_1_1067), 
      .B2(\mem[1] [5]), .ZN(n_1_1_381));
   AOI22_X1 i_1_1_388 (.A1(\mem[92] [5]), .A2(n_1_1_1153), .B1(n_1_1_1108), 
      .B2(\mem[57] [5]), .ZN(n_1_1_382));
   AOI22_X1 i_1_1_389 (.A1(\mem[98] [5]), .A2(n_1_1_1168), .B1(n_1_1_1127), 
      .B2(\mem[72] [5]), .ZN(n_1_1_383));
   AOI22_X1 i_1_1_390 (.A1(\mem[93] [5]), .A2(n_1_1_1155), .B1(n_1_1_1125), 
      .B2(\mem[70] [5]), .ZN(n_1_1_384));
   NOR2_X1 i_1_1_391 (.A1(n_1_1_449), .A2(n_1_1_385), .ZN(n_1_6));
   NOR4_X1 i_1_1_392 (.A1(n_1_1_431), .A2(n_1_1_394), .A3(n_1_1_392), .A4(
      n_1_1_386), .ZN(n_1_1_385));
   NAND4_X1 i_1_1_393 (.A1(n_1_1_428), .A2(n_1_1_424), .A3(n_1_1_391), .A4(
      n_1_1_387), .ZN(n_1_1_386));
   AOI221_X1 i_1_1_394 (.A(n_1_1_388), .B1(n_1_1_1092), .B2(\mem[33] [6]), 
      .C1(\mem[85] [6]), .C2(n_1_1_1058), .ZN(n_1_1_387));
   NAND4_X1 i_1_1_395 (.A1(n_1_1_430), .A2(n_1_1_429), .A3(n_1_1_390), .A4(
      n_1_1_389), .ZN(n_1_1_388));
   AOI22_X1 i_1_1_396 (.A1(\mem[81] [6]), .A2(n_1_1_1139), .B1(n_1_1_1068), 
      .B2(\mem[2] [6]), .ZN(n_1_1_389));
   AOI22_X1 i_1_1_397 (.A1(\mem[49] [6]), .A2(n_1_1_1105), .B1(n_1_1_1030), 
      .B2(\mem[20] [6]), .ZN(n_1_1_390));
   AOI222_X1 i_1_1_398 (.A1(\mem[90] [6]), .A2(n_1_1_1050), .B1(n_1_1_1047), 
      .B2(\mem[83] [6]), .C1(\mem[70] [6]), .C2(n_1_1_1125), .ZN(n_1_1_391));
   NAND4_X1 i_1_1_399 (.A1(n_1_1_423), .A2(n_1_1_422), .A3(n_1_1_418), .A4(
      n_1_1_393), .ZN(n_1_1_392));
   AOI222_X1 i_1_1_400 (.A1(\mem[96] [6]), .A2(n_1_1_1163), .B1(n_1_1_1094), 
      .B2(\mem[35] [6]), .C1(n_1_1_1027), .C2(\mem[27] [6]), .ZN(n_1_1_393));
   NAND4_X1 i_1_1_401 (.A1(n_1_1_427), .A2(n_1_1_417), .A3(n_1_1_399), .A4(
      n_1_1_395), .ZN(n_1_1_394));
   AOI221_X1 i_1_1_402 (.A(n_1_1_396), .B1(n_1_1_1120), .B2(\mem[66] [6]), 
      .C1(\mem[95] [6]), .C2(n_1_1_1053), .ZN(n_1_1_395));
   NAND3_X1 i_1_1_403 (.A1(n_1_1_448), .A2(n_1_1_398), .A3(n_1_1_397), .ZN(
      n_1_1_396));
   AOI22_X1 i_1_1_404 (.A1(\mem[99] [6]), .A2(n_1_1_1171), .B1(n_1_1_1119), 
      .B2(\mem[65] [6]), .ZN(n_1_1_397));
   AOI22_X1 i_1_1_405 (.A1(\mem[11] [6]), .A2(n_1_1_1063), .B1(n_1_1_1062), 
      .B2(\mem[84] [6]), .ZN(n_1_1_398));
   AOI211_X1 i_1_1_406 (.A(n_1_1_410), .B(n_1_1_400), .C1(\mem[8] [6]), .C2(
      n_1_1_1073), .ZN(n_1_1_399));
   NAND3_X1 i_1_1_407 (.A1(read_signal), .A2(n_1_1_406), .A3(n_1_1_401), 
      .ZN(n_1_1_400));
   AOI221_X1 i_1_1_408 (.A(n_1_1_402), .B1(n_1_1_1096), .B2(\mem[37] [6]), 
      .C1(\mem[53] [6]), .C2(n_1_1_1043), .ZN(n_1_1_401));
   NAND3_X1 i_1_1_409 (.A1(n_1_1_405), .A2(n_1_1_404), .A3(n_1_1_403), .ZN(
      n_1_1_402));
   AOI22_X1 i_1_1_410 (.A1(\mem[63] [6]), .A2(n_1_1_1116), .B1(n_1_1_1100), 
      .B2(\mem[41] [6]), .ZN(n_1_1_403));
   AOI22_X1 i_1_1_411 (.A1(\mem[34] [6]), .A2(n_1_1_1093), .B1(n_1_1_1074), 
      .B2(\mem[9] [6]), .ZN(n_1_1_404));
   AOI22_X1 i_1_1_412 (.A1(\mem[13] [6]), .A2(n_1_1_1075), .B1(n_1_1_1032), 
      .B2(\mem[44] [6]), .ZN(n_1_1_405));
   AOI221_X1 i_1_1_413 (.A(n_1_1_407), .B1(n_1_1_1069), .B2(\mem[3] [6]), 
      .C1(\mem[91] [6]), .C2(n_1_1_1037), .ZN(n_1_1_406));
   NAND3_X1 i_1_1_414 (.A1(n_1_1_443), .A2(n_1_1_409), .A3(n_1_1_408), .ZN(
      n_1_1_407));
   AOI22_X1 i_1_1_415 (.A1(\mem[69] [6]), .A2(n_1_1_1123), .B1(n_1_1_1041), 
      .B2(\mem[7] [6]), .ZN(n_1_1_408));
   AOI22_X1 i_1_1_416 (.A1(\mem[68] [6]), .A2(n_1_1_1122), .B1(n_1_1_1042), 
      .B2(\mem[12] [6]), .ZN(n_1_1_409));
   NAND4_X1 i_1_1_417 (.A1(n_1_1_447), .A2(n_1_1_413), .A3(n_1_1_412), .A4(
      n_1_1_411), .ZN(n_1_1_410));
   AOI222_X1 i_1_1_418 (.A1(\mem[72] [6]), .A2(n_1_1_1127), .B1(n_1_1_1104), 
      .B2(\mem[48] [6]), .C1(n_1_1_1097), .C2(\mem[38] [6]), .ZN(n_1_1_411));
   AOI222_X1 i_1_1_419 (.A1(\mem[98] [6]), .A2(n_1_1_1168), .B1(n_1_1_1133), 
      .B2(\mem[77] [6]), .C1(n_1_1_1066), .C2(\mem[0] [6]), .ZN(n_1_1_412));
   AOI221_X1 i_1_1_420 (.A(n_1_1_414), .B1(n_1_1_1142), .B2(\mem[86] [6]), 
      .C1(\mem[97] [6]), .C2(n_1_1_1165), .ZN(n_1_1_413));
   NAND3_X1 i_1_1_421 (.A1(n_1_1_442), .A2(n_1_1_416), .A3(n_1_1_415), .ZN(
      n_1_1_414));
   AOI22_X1 i_1_1_422 (.A1(\mem[73] [6]), .A2(n_1_1_1129), .B1(n_1_1_1055), 
      .B2(\mem[74] [6]), .ZN(n_1_1_415));
   AOI22_X1 i_1_1_423 (.A1(\mem[24] [6]), .A2(n_1_1_1083), .B1(n_1_1_1044), 
      .B2(\mem[26] [6]), .ZN(n_1_1_416));
   AOI22_X1 i_1_1_424 (.A1(\mem[62] [6]), .A2(n_1_1_1029), .B1(n_1_1_1026), 
      .B2(\mem[56] [6]), .ZN(n_1_1_417));
   AOI221_X1 i_1_1_425 (.A(n_1_1_419), .B1(n_1_1_1087), .B2(\mem[30] [6]), 
      .C1(\mem[42] [6]), .C2(n_1_1_1033), .ZN(n_1_1_418));
   NAND3_X1 i_1_1_426 (.A1(n_1_1_445), .A2(n_1_1_421), .A3(n_1_1_420), .ZN(
      n_1_1_419));
   AOI22_X1 i_1_1_427 (.A1(\mem[78] [6]), .A2(n_1_1_1134), .B1(n_1_1_1108), 
      .B2(\mem[57] [6]), .ZN(n_1_1_420));
   AOI22_X1 i_1_1_428 (.A1(\mem[75] [6]), .A2(n_1_1_1061), .B1(n_1_1_1036), 
      .B2(\mem[14] [6]), .ZN(n_1_1_421));
   AOI22_X1 i_1_1_429 (.A1(\mem[80] [6]), .A2(n_1_1_1138), .B1(n_1_1_1101), 
      .B2(\mem[46] [6]), .ZN(n_1_1_422));
   AOI222_X1 i_1_1_430 (.A1(\mem[59] [6]), .A2(n_1_1_1111), .B1(n_1_1_1052), 
      .B2(\mem[23] [6]), .C1(n_1_1_1040), .C2(\mem[52] [6]), .ZN(n_1_1_423));
   AOI221_X1 i_1_1_431 (.A(n_1_1_425), .B1(n_1_1_1088), .B2(\mem[31] [6]), 
      .C1(\mem[51] [6]), .C2(n_1_1_1059), .ZN(n_1_1_424));
   NAND3_X1 i_1_1_432 (.A1(n_1_1_446), .A2(n_1_1_444), .A3(n_1_1_426), .ZN(
      n_1_1_425));
   AOI22_X1 i_1_1_433 (.A1(\mem[25] [6]), .A2(n_1_1_1084), .B1(n_1_1_1038), 
      .B2(\mem[15] [6]), .ZN(n_1_1_426));
   AOI22_X1 i_1_1_434 (.A1(\mem[87] [6]), .A2(n_1_1_1144), .B1(n_1_1_1035), 
      .B2(\mem[50] [6]), .ZN(n_1_1_427));
   AOI222_X1 i_1_1_435 (.A1(\mem[79] [6]), .A2(n_1_1_1135), .B1(n_1_1_1051), 
      .B2(\mem[29] [6]), .C1(n_1_1_1028), .C2(\mem[82] [6]), .ZN(n_1_1_428));
   AOI22_X1 i_1_1_436 (.A1(\mem[6] [6]), .A2(n_1_1_1072), .B1(n_1_1_1071), 
      .B2(\mem[5] [6]), .ZN(n_1_1_429));
   AOI22_X1 i_1_1_437 (.A1(\mem[36] [6]), .A2(n_1_1_1095), .B1(n_1_1_1048), 
      .B2(\mem[10] [6]), .ZN(n_1_1_430));
   NAND2_X1 i_1_1_438 (.A1(n_1_1_437), .A2(n_1_1_432), .ZN(n_1_1_431));
   AOI221_X1 i_1_1_439 (.A(n_1_1_433), .B1(n_1_1_1106), .B2(\mem[54] [6]), 
      .C1(\mem[89] [6]), .C2(n_1_1_1148), .ZN(n_1_1_432));
   NAND3_X1 i_1_1_440 (.A1(n_1_1_436), .A2(n_1_1_435), .A3(n_1_1_434), .ZN(
      n_1_1_433));
   AOI22_X1 i_1_1_441 (.A1(\mem[94] [6]), .A2(n_1_1_1157), .B1(n_1_1_1049), 
      .B2(\mem[17] [6]), .ZN(n_1_1_434));
   AOI22_X1 i_1_1_442 (.A1(\mem[100] [6]), .A2(n_1_1_1174), .B1(n_1_1_1039), 
      .B2(\mem[76] [6]), .ZN(n_1_1_435));
   AOI22_X1 i_1_1_443 (.A1(\mem[55] [6]), .A2(n_1_1_1107), .B1(n_1_1_1091), 
      .B2(\mem[32] [6]), .ZN(n_1_1_436));
   AOI221_X1 i_1_1_444 (.A(n_1_1_438), .B1(n_1_1_1080), .B2(\mem[19] [6]), 
      .C1(\mem[93] [6]), .C2(n_1_1_1155), .ZN(n_1_1_437));
   NAND3_X1 i_1_1_445 (.A1(n_1_1_441), .A2(n_1_1_440), .A3(n_1_1_439), .ZN(
      n_1_1_438));
   AOI22_X1 i_1_1_446 (.A1(\mem[28] [6]), .A2(n_1_1_1060), .B1(n_1_1_1054), 
      .B2(\mem[22] [6]), .ZN(n_1_1_439));
   AOI22_X1 i_1_1_447 (.A1(\mem[92] [6]), .A2(n_1_1_1153), .B1(n_1_1_1064), 
      .B2(\mem[18] [6]), .ZN(n_1_1_440));
   AOI22_X1 i_1_1_448 (.A1(\mem[71] [6]), .A2(n_1_1_1126), .B1(n_1_1_1109), 
      .B2(\mem[58] [6]), .ZN(n_1_1_441));
   AOI22_X1 i_1_1_449 (.A1(\mem[21] [6]), .A2(n_1_1_1081), .B1(n_1_1_1046), 
      .B2(\mem[60] [6]), .ZN(n_1_1_442));
   AOI22_X1 i_1_1_450 (.A1(\mem[45] [6]), .A2(n_1_1_1045), .B1(n_1_1_1025), 
      .B2(\mem[43] [6]), .ZN(n_1_1_443));
   AOI22_X1 i_1_1_451 (.A1(\mem[67] [6]), .A2(n_1_1_1121), .B1(n_1_1_1031), 
      .B2(\mem[39] [6]), .ZN(n_1_1_444));
   AOI22_X1 i_1_1_452 (.A1(\mem[1] [6]), .A2(n_1_1_1067), .B1(n_1_1_1056), 
      .B2(\mem[88] [6]), .ZN(n_1_1_445));
   AOI22_X1 i_1_1_453 (.A1(\mem[47] [6]), .A2(n_1_1_1102), .B1(n_1_1_1078), 
      .B2(\mem[16] [6]), .ZN(n_1_1_446));
   AOI22_X1 i_1_1_454 (.A1(\mem[40] [6]), .A2(n_1_1_1099), .B1(n_1_1_1057), 
      .B2(\mem[61] [6]), .ZN(n_1_1_447));
   AOI22_X1 i_1_1_455 (.A1(\mem[64] [6]), .A2(n_1_1_1118), .B1(n_1_1_1070), 
      .B2(\mem[4] [6]), .ZN(n_1_1_448));
   NOR2_X1 i_1_1_456 (.A1(read_signal), .A2(dataout[6]), .ZN(n_1_1_449));
   AOI21_X1 i_1_1_457 (.A(n_1_1_513), .B1(n_1_1_501), .B2(n_1_1_450), .ZN(n_1_7));
   NOR4_X1 i_1_1_458 (.A1(n_1_1_497), .A2(n_1_1_480), .A3(n_1_1_466), .A4(
      n_1_1_451), .ZN(n_1_1_450));
   NAND4_X1 i_1_1_459 (.A1(n_1_1_507), .A2(n_1_1_465), .A3(n_1_1_460), .A4(
      n_1_1_452), .ZN(n_1_1_451));
   AOI221_X1 i_1_1_460 (.A(n_1_1_453), .B1(n_1_1_1030), .B2(\mem[20] [7]), 
      .C1(\mem[60] [7]), .C2(n_1_1_1046), .ZN(n_1_1_452));
   NAND3_X1 i_1_1_461 (.A1(read_signal), .A2(n_1_1_506), .A3(n_1_1_454), 
      .ZN(n_1_1_453));
   AOI21_X1 i_1_1_462 (.A(n_1_1_455), .B1(n_1_1_1105), .B2(\mem[49] [7]), 
      .ZN(n_1_1_454));
   NAND4_X1 i_1_1_463 (.A1(n_1_1_459), .A2(n_1_1_458), .A3(n_1_1_457), .A4(
      n_1_1_456), .ZN(n_1_1_455));
   AOI22_X1 i_1_1_464 (.A1(\mem[16] [7]), .A2(n_1_1_1078), .B1(n_1_1_1057), 
      .B2(\mem[61] [7]), .ZN(n_1_1_456));
   AOI22_X1 i_1_1_465 (.A1(\mem[36] [7]), .A2(n_1_1_1095), .B1(n_1_1_1058), 
      .B2(\mem[85] [7]), .ZN(n_1_1_457));
   AOI22_X1 i_1_1_466 (.A1(\mem[77] [7]), .A2(n_1_1_1133), .B1(n_1_1_1099), 
      .B2(\mem[40] [7]), .ZN(n_1_1_458));
   AOI22_X1 i_1_1_467 (.A1(\mem[79] [7]), .A2(n_1_1_1135), .B1(n_1_1_1052), 
      .B2(\mem[23] [7]), .ZN(n_1_1_459));
   AOI221_X1 i_1_1_468 (.A(n_1_1_461), .B1(n_1_1_1063), .B2(\mem[11] [7]), 
      .C1(\mem[44] [7]), .C2(n_1_1_1032), .ZN(n_1_1_460));
   NAND3_X1 i_1_1_469 (.A1(n_1_1_464), .A2(n_1_1_463), .A3(n_1_1_462), .ZN(
      n_1_1_461));
   AOI222_X1 i_1_1_470 (.A1(\mem[97] [7]), .A2(n_1_1_1165), .B1(n_1_1_1111), 
      .B2(\mem[59] [7]), .C1(n_1_1_1029), .C2(\mem[62] [7]), .ZN(n_1_1_462));
   AOI22_X1 i_1_1_471 (.A1(\mem[75] [7]), .A2(n_1_1_1061), .B1(n_1_1_1040), 
      .B2(\mem[52] [7]), .ZN(n_1_1_463));
   AOI222_X1 i_1_1_472 (.A1(\mem[65] [7]), .A2(n_1_1_1119), .B1(n_1_1_1101), 
      .B2(\mem[46] [7]), .C1(n_1_1_1100), .C2(\mem[41] [7]), .ZN(n_1_1_464));
   AOI222_X1 i_1_1_473 (.A1(\mem[78] [7]), .A2(n_1_1_1134), .B1(n_1_1_1026), 
      .B2(\mem[56] [7]), .C1(n_1_1_1037), .C2(\mem[91] [7]), .ZN(n_1_1_465));
   NAND4_X1 i_1_1_474 (.A1(n_1_1_479), .A2(n_1_1_478), .A3(n_1_1_473), .A4(
      n_1_1_467), .ZN(n_1_1_466));
   AOI221_X1 i_1_1_475 (.A(n_1_1_468), .B1(n_1_1_1044), .B2(\mem[26] [7]), 
      .C1(\mem[70] [7]), .C2(n_1_1_1125), .ZN(n_1_1_467));
   NAND4_X1 i_1_1_476 (.A1(n_1_1_472), .A2(n_1_1_471), .A3(n_1_1_470), .A4(
      n_1_1_469), .ZN(n_1_1_468));
   AOI22_X1 i_1_1_477 (.A1(\mem[24] [7]), .A2(n_1_1_1083), .B1(n_1_1_1036), 
      .B2(\mem[14] [7]), .ZN(n_1_1_469));
   AOI22_X1 i_1_1_478 (.A1(\mem[72] [7]), .A2(n_1_1_1127), .B1(n_1_1_1080), 
      .B2(\mem[19] [7]), .ZN(n_1_1_470));
   AOI22_X1 i_1_1_479 (.A1(\mem[18] [7]), .A2(n_1_1_1064), .B1(n_1_1_1039), 
      .B2(\mem[76] [7]), .ZN(n_1_1_471));
   AOI22_X1 i_1_1_480 (.A1(\mem[81] [7]), .A2(n_1_1_1139), .B1(n_1_1_1049), 
      .B2(\mem[17] [7]), .ZN(n_1_1_472));
   AOI221_X1 i_1_1_481 (.A(n_1_1_474), .B1(n_1_1_1096), .B2(\mem[37] [7]), 
      .C1(\mem[45] [7]), .C2(n_1_1_1045), .ZN(n_1_1_473));
   NAND3_X1 i_1_1_482 (.A1(n_1_1_477), .A2(n_1_1_476), .A3(n_1_1_475), .ZN(
      n_1_1_474));
   AOI22_X1 i_1_1_483 (.A1(\mem[53] [7]), .A2(n_1_1_1043), .B1(n_1_1_1031), 
      .B2(\mem[39] [7]), .ZN(n_1_1_475));
   AOI22_X1 i_1_1_484 (.A1(\mem[35] [7]), .A2(n_1_1_1094), .B1(n_1_1_1074), 
      .B2(\mem[9] [7]), .ZN(n_1_1_476));
   AOI22_X1 i_1_1_485 (.A1(\mem[68] [7]), .A2(n_1_1_1122), .B1(n_1_1_1059), 
      .B2(\mem[51] [7]), .ZN(n_1_1_477));
   AOI222_X1 i_1_1_486 (.A1(\mem[73] [7]), .A2(n_1_1_1129), .B1(n_1_1_1087), 
      .B2(\mem[30] [7]), .C1(n_1_1_1073), .C2(\mem[8] [7]), .ZN(n_1_1_478));
   AOI222_X1 i_1_1_487 (.A1(\mem[80] [7]), .A2(n_1_1_1138), .B1(n_1_1_1066), 
      .B2(\mem[0] [7]), .C1(n_1_1_1055), .C2(\mem[74] [7]), .ZN(n_1_1_479));
   NAND4_X1 i_1_1_488 (.A1(n_1_1_492), .A2(n_1_1_487), .A3(n_1_1_484), .A4(
      n_1_1_481), .ZN(n_1_1_480));
   AOI221_X1 i_1_1_489 (.A(n_1_1_482), .B1(n_1_1_1048), .B2(\mem[10] [7]), 
      .C1(\mem[82] [7]), .C2(n_1_1_1028), .ZN(n_1_1_481));
   NAND3_X1 i_1_1_490 (.A1(n_1_1_510), .A2(n_1_1_509), .A3(n_1_1_483), .ZN(
      n_1_1_482));
   AOI22_X1 i_1_1_491 (.A1(\mem[93] [7]), .A2(n_1_1_1155), .B1(n_1_1_1123), 
      .B2(\mem[69] [7]), .ZN(n_1_1_483));
   AOI221_X1 i_1_1_492 (.A(n_1_1_485), .B1(n_1_1_1107), .B2(\mem[55] [7]), 
      .C1(\mem[58] [7]), .C2(n_1_1_1109), .ZN(n_1_1_484));
   NAND3_X1 i_1_1_493 (.A1(n_1_1_511), .A2(n_1_1_508), .A3(n_1_1_486), .ZN(
      n_1_1_485));
   AOI22_X1 i_1_1_494 (.A1(\mem[25] [7]), .A2(n_1_1_1084), .B1(n_1_1_1067), 
      .B2(\mem[1] [7]), .ZN(n_1_1_486));
   AOI221_X1 i_1_1_495 (.A(n_1_1_488), .B1(n_1_1_1070), .B2(\mem[4] [7]), 
      .C1(\mem[67] [7]), .C2(n_1_1_1121), .ZN(n_1_1_487));
   NAND3_X1 i_1_1_496 (.A1(n_1_1_491), .A2(n_1_1_490), .A3(n_1_1_489), .ZN(
      n_1_1_488));
   AOI22_X1 i_1_1_497 (.A1(\mem[66] [7]), .A2(n_1_1_1120), .B1(n_1_1_1053), 
      .B2(\mem[95] [7]), .ZN(n_1_1_489));
   AOI22_X1 i_1_1_498 (.A1(\mem[96] [7]), .A2(n_1_1_1163), .B1(n_1_1_1081), 
      .B2(\mem[21] [7]), .ZN(n_1_1_490));
   AOI22_X1 i_1_1_499 (.A1(\mem[99] [7]), .A2(n_1_1_1171), .B1(n_1_1_1069), 
      .B2(\mem[3] [7]), .ZN(n_1_1_491));
   AOI221_X1 i_1_1_500 (.A(n_1_1_493), .B1(n_1_1_1126), .B2(\mem[71] [7]), 
      .C1(\mem[90] [7]), .C2(n_1_1_1050), .ZN(n_1_1_492));
   NAND3_X1 i_1_1_501 (.A1(n_1_1_496), .A2(n_1_1_495), .A3(n_1_1_494), .ZN(
      n_1_1_493));
   AOI22_X1 i_1_1_502 (.A1(\mem[33] [7]), .A2(n_1_1_1092), .B1(n_1_1_1051), 
      .B2(\mem[29] [7]), .ZN(n_1_1_494));
   AOI22_X1 i_1_1_503 (.A1(\mem[87] [7]), .A2(n_1_1_1144), .B1(n_1_1_1062), 
      .B2(\mem[84] [7]), .ZN(n_1_1_495));
   AOI22_X1 i_1_1_504 (.A1(\mem[83] [7]), .A2(n_1_1_1047), .B1(n_1_1_1042), 
      .B2(\mem[12] [7]), .ZN(n_1_1_496));
   NAND4_X1 i_1_1_505 (.A1(n_1_1_512), .A2(n_1_1_500), .A3(n_1_1_499), .A4(
      n_1_1_498), .ZN(n_1_1_497));
   AOI22_X1 i_1_1_506 (.A1(\mem[47] [7]), .A2(n_1_1_1102), .B1(n_1_1_1075), 
      .B2(\mem[13] [7]), .ZN(n_1_1_498));
   AOI22_X1 i_1_1_507 (.A1(\mem[63] [7]), .A2(n_1_1_1116), .B1(n_1_1_1088), 
      .B2(\mem[31] [7]), .ZN(n_1_1_499));
   AOI22_X1 i_1_1_508 (.A1(\mem[54] [7]), .A2(n_1_1_1106), .B1(n_1_1_1033), 
      .B2(\mem[42] [7]), .ZN(n_1_1_500));
   AOI221_X1 i_1_1_509 (.A(n_1_1_502), .B1(n_1_1_1093), .B2(\mem[34] [7]), 
      .C1(\mem[38] [7]), .C2(n_1_1_1097), .ZN(n_1_1_501));
   NAND3_X1 i_1_1_510 (.A1(n_1_1_505), .A2(n_1_1_504), .A3(n_1_1_503), .ZN(
      n_1_1_502));
   AOI22_X1 i_1_1_511 (.A1(\mem[100] [7]), .A2(n_1_1_1174), .B1(n_1_1_1035), 
      .B2(\mem[50] [7]), .ZN(n_1_1_503));
   AOI22_X1 i_1_1_512 (.A1(\mem[48] [7]), .A2(n_1_1_1104), .B1(n_1_1_1025), 
      .B2(\mem[43] [7]), .ZN(n_1_1_504));
   AOI22_X1 i_1_1_513 (.A1(\mem[98] [7]), .A2(n_1_1_1168), .B1(n_1_1_1068), 
      .B2(\mem[2] [7]), .ZN(n_1_1_505));
   AOI22_X1 i_1_1_514 (.A1(\mem[92] [7]), .A2(n_1_1_1153), .B1(n_1_1_1091), 
      .B2(\mem[32] [7]), .ZN(n_1_1_506));
   AOI222_X1 i_1_1_515 (.A1(\mem[94] [7]), .A2(n_1_1_1157), .B1(n_1_1_1054), 
      .B2(\mem[22] [7]), .C1(n_1_1_1038), .C2(\mem[15] [7]), .ZN(n_1_1_507));
   AOI22_X1 i_1_1_516 (.A1(\mem[57] [7]), .A2(n_1_1_1108), .B1(n_1_1_1027), 
      .B2(\mem[27] [7]), .ZN(n_1_1_508));
   AOI22_X1 i_1_1_517 (.A1(\mem[89] [7]), .A2(n_1_1_1148), .B1(n_1_1_1056), 
      .B2(\mem[88] [7]), .ZN(n_1_1_509));
   AOI22_X1 i_1_1_518 (.A1(\mem[86] [7]), .A2(n_1_1_1142), .B1(n_1_1_1072), 
      .B2(\mem[6] [7]), .ZN(n_1_1_510));
   AOI22_X1 i_1_1_519 (.A1(\mem[5] [7]), .A2(n_1_1_1071), .B1(n_1_1_1041), 
      .B2(\mem[7] [7]), .ZN(n_1_1_511));
   AOI22_X1 i_1_1_520 (.A1(\mem[64] [7]), .A2(n_1_1_1118), .B1(n_1_1_1060), 
      .B2(\mem[28] [7]), .ZN(n_1_1_512));
   NOR2_X1 i_1_1_521 (.A1(read_signal), .A2(dataout[7]), .ZN(n_1_1_513));
   MUX2_X1 i_1_1_522 (.A(dataout[8]), .B(n_1_1_514), .S(read_signal), .Z(n_1_8));
   NAND4_X1 i_1_1_523 (.A1(n_1_1_561), .A2(n_1_1_532), .A3(n_1_1_520), .A4(
      n_1_1_515), .ZN(n_1_1_514));
   AOI221_X1 i_1_1_524 (.A(n_1_1_516), .B1(n_1_1_1066), .B2(\mem[0] [8]), 
      .C1(\mem[89] [8]), .C2(n_1_1_1148), .ZN(n_1_1_515));
   NAND3_X1 i_1_1_525 (.A1(n_1_1_519), .A2(n_1_1_518), .A3(n_1_1_517), .ZN(
      n_1_1_516));
   AOI22_X1 i_1_1_526 (.A1(\mem[99] [8]), .A2(n_1_1_1171), .B1(n_1_1_1056), 
      .B2(\mem[88] [8]), .ZN(n_1_1_517));
   AOI22_X1 i_1_1_527 (.A1(\mem[98] [8]), .A2(n_1_1_1168), .B1(n_1_1_1093), 
      .B2(\mem[34] [8]), .ZN(n_1_1_518));
   AOI22_X1 i_1_1_528 (.A1(\mem[92] [8]), .A2(n_1_1_1153), .B1(n_1_1_1051), 
      .B2(\mem[29] [8]), .ZN(n_1_1_519));
   AOI221_X1 i_1_1_529 (.A(n_1_1_521), .B1(n_1_1_1078), .B2(\mem[16] [8]), 
      .C1(\mem[84] [8]), .C2(n_1_1_1062), .ZN(n_1_1_520));
   NAND4_X1 i_1_1_530 (.A1(n_1_1_530), .A2(n_1_1_529), .A3(n_1_1_528), .A4(
      n_1_1_522), .ZN(n_1_1_521));
   AOI221_X1 i_1_1_531 (.A(n_1_1_523), .B1(n_1_1_1052), .B2(\mem[23] [8]), 
      .C1(\mem[75] [8]), .C2(n_1_1_1061), .ZN(n_1_1_522));
   NAND4_X1 i_1_1_532 (.A1(n_1_1_527), .A2(n_1_1_526), .A3(n_1_1_525), .A4(
      n_1_1_524), .ZN(n_1_1_523));
   AOI22_X1 i_1_1_533 (.A1(\mem[31] [8]), .A2(n_1_1_1088), .B1(n_1_1_1041), 
      .B2(\mem[7] [8]), .ZN(n_1_1_524));
   AOI22_X1 i_1_1_534 (.A1(\mem[79] [8]), .A2(n_1_1_1135), .B1(n_1_1_1071), 
      .B2(\mem[5] [8]), .ZN(n_1_1_525));
   AOI22_X1 i_1_1_535 (.A1(\mem[2] [8]), .A2(n_1_1_1068), .B1(n_1_1_1058), 
      .B2(\mem[85] [8]), .ZN(n_1_1_526));
   AOI22_X1 i_1_1_536 (.A1(\mem[32] [8]), .A2(n_1_1_1091), .B1(n_1_1_1030), 
      .B2(\mem[20] [8]), .ZN(n_1_1_527));
   AOI22_X1 i_1_1_537 (.A1(\mem[35] [8]), .A2(n_1_1_1094), .B1(n_1_1_1026), 
      .B2(\mem[56] [8]), .ZN(n_1_1_528));
   AOI222_X1 i_1_1_538 (.A1(\mem[67] [8]), .A2(n_1_1_1121), .B1(n_1_1_1116), 
      .B2(\mem[63] [8]), .C1(n_1_1_1038), .C2(\mem[15] [8]), .ZN(n_1_1_529));
   AOI221_X1 i_1_1_539 (.A(n_1_1_531), .B1(n_1_1_1100), .B2(\mem[41] [8]), 
      .C1(\mem[95] [8]), .C2(n_1_1_1053), .ZN(n_1_1_530));
   NAND4_X1 i_1_1_540 (.A1(n_1_1_573), .A2(n_1_1_568), .A3(n_1_1_560), .A4(
      n_1_1_558), .ZN(n_1_1_531));
   NOR3_X1 i_1_1_541 (.A1(n_1_1_555), .A2(n_1_1_534), .A3(n_1_1_533), .ZN(
      n_1_1_532));
   NAND4_X1 i_1_1_542 (.A1(n_1_1_572), .A2(n_1_1_569), .A3(n_1_1_562), .A4(
      n_1_1_559), .ZN(n_1_1_533));
   NAND4_X1 i_1_1_543 (.A1(n_1_1_554), .A2(n_1_1_548), .A3(n_1_1_547), .A4(
      n_1_1_535), .ZN(n_1_1_534));
   NOR3_X1 i_1_1_544 (.A1(n_1_1_538), .A2(n_1_1_537), .A3(n_1_1_536), .ZN(
      n_1_1_535));
   NAND4_X1 i_1_1_545 (.A1(n_1_1_575), .A2(n_1_1_574), .A3(n_1_1_571), .A4(
      n_1_1_556), .ZN(n_1_1_536));
   NAND4_X1 i_1_1_546 (.A1(n_1_1_576), .A2(n_1_1_567), .A3(n_1_1_566), .A4(
      n_1_1_557), .ZN(n_1_1_537));
   NAND4_X1 i_1_1_547 (.A1(n_1_1_546), .A2(n_1_1_545), .A3(n_1_1_540), .A4(
      n_1_1_539), .ZN(n_1_1_538));
   AOI222_X1 i_1_1_548 (.A1(\mem[58] [8]), .A2(n_1_1_1109), .B1(n_1_1_1070), 
      .B2(\mem[4] [8]), .C1(n_1_1_1049), .C2(\mem[17] [8]), .ZN(n_1_1_539));
   AOI221_X1 i_1_1_549 (.A(n_1_1_541), .B1(n_1_1_1059), .B2(\mem[51] [8]), 
      .C1(\mem[52] [8]), .C2(n_1_1_1040), .ZN(n_1_1_540));
   NAND3_X1 i_1_1_550 (.A1(n_1_1_544), .A2(n_1_1_543), .A3(n_1_1_542), .ZN(
      n_1_1_541));
   AOI22_X1 i_1_1_551 (.A1(\mem[38] [8]), .A2(n_1_1_1097), .B1(n_1_1_1072), 
      .B2(\mem[6] [8]), .ZN(n_1_1_542));
   AOI22_X1 i_1_1_552 (.A1(\mem[57] [8]), .A2(n_1_1_1108), .B1(n_1_1_1101), 
      .B2(\mem[46] [8]), .ZN(n_1_1_543));
   AOI22_X1 i_1_1_553 (.A1(\mem[25] [8]), .A2(n_1_1_1084), .B1(n_1_1_1063), 
      .B2(\mem[11] [8]), .ZN(n_1_1_544));
   AOI22_X1 i_1_1_554 (.A1(\mem[66] [8]), .A2(n_1_1_1120), .B1(n_1_1_1037), 
      .B2(\mem[91] [8]), .ZN(n_1_1_545));
   AOI222_X1 i_1_1_555 (.A1(\mem[24] [8]), .A2(n_1_1_1083), .B1(n_1_1_1069), 
      .B2(\mem[3] [8]), .C1(n_1_1_1067), .C2(\mem[1] [8]), .ZN(n_1_1_546));
   AOI222_X1 i_1_1_556 (.A1(\mem[22] [8]), .A2(n_1_1_1054), .B1(n_1_1_1036), 
      .B2(\mem[14] [8]), .C1(n_1_1_1045), .C2(\mem[45] [8]), .ZN(n_1_1_547));
   AOI221_X1 i_1_1_557 (.A(n_1_1_549), .B1(n_1_1_1157), .B2(\mem[94] [8]), 
      .C1(\mem[97] [8]), .C2(n_1_1_1165), .ZN(n_1_1_548));
   NAND4_X1 i_1_1_558 (.A1(n_1_1_553), .A2(n_1_1_552), .A3(n_1_1_551), .A4(
      n_1_1_550), .ZN(n_1_1_549));
   AOI22_X1 i_1_1_559 (.A1(\mem[73] [8]), .A2(n_1_1_1129), .B1(n_1_1_1031), 
      .B2(\mem[39] [8]), .ZN(n_1_1_550));
   AOI22_X1 i_1_1_560 (.A1(\mem[60] [8]), .A2(n_1_1_1046), .B1(n_1_1_1039), 
      .B2(\mem[76] [8]), .ZN(n_1_1_551));
   AOI22_X1 i_1_1_561 (.A1(\mem[30] [8]), .A2(n_1_1_1087), .B1(n_1_1_1047), 
      .B2(\mem[83] [8]), .ZN(n_1_1_552));
   AOI22_X1 i_1_1_562 (.A1(\mem[81] [8]), .A2(n_1_1_1139), .B1(n_1_1_1126), 
      .B2(\mem[71] [8]), .ZN(n_1_1_553));
   AOI222_X1 i_1_1_563 (.A1(\mem[69] [8]), .A2(n_1_1_1123), .B1(n_1_1_1035), 
      .B2(\mem[50] [8]), .C1(n_1_1_1025), .C2(\mem[43] [8]), .ZN(n_1_1_554));
   NAND4_X1 i_1_1_564 (.A1(n_1_1_570), .A2(n_1_1_565), .A3(n_1_1_564), .A4(
      n_1_1_563), .ZN(n_1_1_555));
   AOI22_X1 i_1_1_565 (.A1(\mem[80] [8]), .A2(n_1_1_1138), .B1(n_1_1_1048), 
      .B2(\mem[10] [8]), .ZN(n_1_1_556));
   AOI22_X1 i_1_1_566 (.A1(\mem[54] [8]), .A2(n_1_1_1106), .B1(n_1_1_1027), 
      .B2(\mem[27] [8]), .ZN(n_1_1_557));
   AOI22_X1 i_1_1_567 (.A1(\mem[96] [8]), .A2(n_1_1_1163), .B1(n_1_1_1155), 
      .B2(\mem[93] [8]), .ZN(n_1_1_558));
   AOI22_X1 i_1_1_568 (.A1(\mem[68] [8]), .A2(n_1_1_1122), .B1(n_1_1_1075), 
      .B2(\mem[13] [8]), .ZN(n_1_1_559));
   AOI22_X1 i_1_1_569 (.A1(\mem[64] [8]), .A2(n_1_1_1118), .B1(n_1_1_1057), 
      .B2(\mem[61] [8]), .ZN(n_1_1_560));
   AOI22_X1 i_1_1_570 (.A1(\mem[87] [8]), .A2(n_1_1_1144), .B1(n_1_1_1134), 
      .B2(\mem[78] [8]), .ZN(n_1_1_561));
   AOI22_X1 i_1_1_571 (.A1(\mem[55] [8]), .A2(n_1_1_1107), .B1(n_1_1_1064), 
      .B2(\mem[18] [8]), .ZN(n_1_1_562));
   AOI22_X1 i_1_1_572 (.A1(\mem[59] [8]), .A2(n_1_1_1111), .B1(n_1_1_1074), 
      .B2(\mem[9] [8]), .ZN(n_1_1_563));
   AOI22_X1 i_1_1_573 (.A1(\mem[37] [8]), .A2(n_1_1_1096), .B1(n_1_1_1080), 
      .B2(\mem[19] [8]), .ZN(n_1_1_564));
   AOI22_X1 i_1_1_574 (.A1(\mem[47] [8]), .A2(n_1_1_1102), .B1(n_1_1_1081), 
      .B2(\mem[21] [8]), .ZN(n_1_1_565));
   AOI22_X1 i_1_1_575 (.A1(\mem[77] [8]), .A2(n_1_1_1133), .B1(n_1_1_1104), 
      .B2(\mem[48] [8]), .ZN(n_1_1_566));
   AOI22_X1 i_1_1_576 (.A1(\mem[8] [8]), .A2(n_1_1_1073), .B1(n_1_1_1033), 
      .B2(\mem[42] [8]), .ZN(n_1_1_567));
   AOI22_X1 i_1_1_577 (.A1(\mem[72] [8]), .A2(n_1_1_1127), .B1(n_1_1_1044), 
      .B2(\mem[26] [8]), .ZN(n_1_1_568));
   AOI22_X1 i_1_1_578 (.A1(\mem[53] [8]), .A2(n_1_1_1043), .B1(n_1_1_1032), 
      .B2(\mem[44] [8]), .ZN(n_1_1_569));
   AOI22_X1 i_1_1_579 (.A1(\mem[40] [8]), .A2(n_1_1_1099), .B1(n_1_1_1095), 
      .B2(\mem[36] [8]), .ZN(n_1_1_570));
   AOI22_X1 i_1_1_580 (.A1(\mem[90] [8]), .A2(n_1_1_1050), .B1(n_1_1_1042), 
      .B2(\mem[12] [8]), .ZN(n_1_1_571));
   AOI22_X1 i_1_1_581 (.A1(\mem[70] [8]), .A2(n_1_1_1125), .B1(n_1_1_1060), 
      .B2(\mem[28] [8]), .ZN(n_1_1_572));
   AOI22_X1 i_1_1_582 (.A1(\mem[49] [8]), .A2(n_1_1_1105), .B1(n_1_1_1028), 
      .B2(\mem[82] [8]), .ZN(n_1_1_573));
   AOI22_X1 i_1_1_583 (.A1(\mem[100] [8]), .A2(n_1_1_1174), .B1(n_1_1_1092), 
      .B2(\mem[33] [8]), .ZN(n_1_1_574));
   AOI22_X1 i_1_1_584 (.A1(\mem[86] [8]), .A2(n_1_1_1142), .B1(n_1_1_1055), 
      .B2(\mem[74] [8]), .ZN(n_1_1_575));
   AOI22_X1 i_1_1_585 (.A1(\mem[65] [8]), .A2(n_1_1_1119), .B1(n_1_1_1029), 
      .B2(\mem[62] [8]), .ZN(n_1_1_576));
   INV_X1 i_1_1_586 (.A(n_1_1_577), .ZN(n_1_9));
   OAI22_X1 i_1_1_587 (.A1(n_1_1_584), .A2(n_1_1_578), .B1(read_signal), 
      .B2(dataout[9]), .ZN(n_1_1_577));
   NAND4_X1 i_1_1_588 (.A1(n_1_1_638), .A2(n_1_1_628), .A3(n_1_1_580), .A4(
      n_1_1_579), .ZN(n_1_1_578));
   AOI222_X1 i_1_1_589 (.A1(\mem[96] [9]), .A2(n_1_1_1163), .B1(n_1_1_1139), 
      .B2(\mem[81] [9]), .C1(n_1_1_1054), .C2(\mem[22] [9]), .ZN(n_1_1_579));
   AOI221_X1 i_1_1_590 (.A(n_1_1_581), .B1(n_1_1_1084), .B2(\mem[25] [9]), 
      .C1(\mem[79] [9]), .C2(n_1_1_1135), .ZN(n_1_1_580));
   NAND3_X1 i_1_1_591 (.A1(n_1_1_637), .A2(n_1_1_583), .A3(n_1_1_582), .ZN(
      n_1_1_581));
   AOI222_X1 i_1_1_592 (.A1(\mem[94] [9]), .A2(n_1_1_1157), .B1(n_1_1_1138), 
      .B2(\mem[80] [9]), .C1(n_1_1_1093), .C2(\mem[34] [9]), .ZN(n_1_1_582));
   AOI222_X1 i_1_1_593 (.A1(\mem[99] [9]), .A2(n_1_1_1171), .B1(n_1_1_1073), 
      .B2(\mem[8] [9]), .C1(n_1_1_1056), .C2(\mem[88] [9]), .ZN(n_1_1_583));
   NAND3_X1 i_1_1_594 (.A1(n_1_1_632), .A2(n_1_1_604), .A3(n_1_1_585), .ZN(
      n_1_1_584));
   AND4_X1 i_1_1_595 (.A1(n_1_1_599), .A2(n_1_1_593), .A3(n_1_1_587), .A4(
      n_1_1_586), .ZN(n_1_1_585));
   AOI222_X1 i_1_1_596 (.A1(\mem[64] [9]), .A2(n_1_1_1118), .B1(n_1_1_1067), 
      .B2(\mem[1] [9]), .C1(n_1_1_1043), .C2(\mem[53] [9]), .ZN(n_1_1_586));
   AOI221_X1 i_1_1_597 (.A(n_1_1_588), .B1(n_1_1_1107), .B2(\mem[55] [9]), 
      .C1(\mem[60] [9]), .C2(n_1_1_1046), .ZN(n_1_1_587));
   NAND4_X1 i_1_1_598 (.A1(n_1_1_592), .A2(n_1_1_591), .A3(n_1_1_590), .A4(
      n_1_1_589), .ZN(n_1_1_588));
   AOI22_X1 i_1_1_599 (.A1(\mem[100] [9]), .A2(n_1_1_1174), .B1(n_1_1_1127), 
      .B2(\mem[72] [9]), .ZN(n_1_1_589));
   AOI22_X1 i_1_1_600 (.A1(\mem[87] [9]), .A2(n_1_1_1144), .B1(n_1_1_1105), 
      .B2(\mem[49] [9]), .ZN(n_1_1_590));
   AOI22_X1 i_1_1_601 (.A1(\mem[6] [9]), .A2(n_1_1_1072), .B1(n_1_1_1047), 
      .B2(\mem[83] [9]), .ZN(n_1_1_591));
   AOI22_X1 i_1_1_602 (.A1(\mem[70] [9]), .A2(n_1_1_1125), .B1(n_1_1_1040), 
      .B2(\mem[52] [9]), .ZN(n_1_1_592));
   AOI221_X1 i_1_1_603 (.A(n_1_1_594), .B1(n_1_1_1116), .B2(\mem[63] [9]), 
      .C1(\mem[73] [9]), .C2(n_1_1_1129), .ZN(n_1_1_593));
   NAND4_X1 i_1_1_604 (.A1(n_1_1_598), .A2(n_1_1_597), .A3(n_1_1_596), .A4(
      n_1_1_595), .ZN(n_1_1_594));
   AOI22_X1 i_1_1_605 (.A1(\mem[41] [9]), .A2(n_1_1_1100), .B1(n_1_1_1030), 
      .B2(\mem[20] [9]), .ZN(n_1_1_595));
   AOI22_X1 i_1_1_606 (.A1(\mem[68] [9]), .A2(n_1_1_1122), .B1(n_1_1_1074), 
      .B2(\mem[9] [9]), .ZN(n_1_1_596));
   AOI22_X1 i_1_1_607 (.A1(\mem[21] [9]), .A2(n_1_1_1081), .B1(n_1_1_1057), 
      .B2(\mem[61] [9]), .ZN(n_1_1_597));
   AOI22_X1 i_1_1_608 (.A1(\mem[59] [9]), .A2(n_1_1_1111), .B1(n_1_1_1088), 
      .B2(\mem[31] [9]), .ZN(n_1_1_598));
   AOI221_X1 i_1_1_609 (.A(n_1_1_600), .B1(n_1_1_1075), .B2(\mem[13] [9]), 
      .C1(\mem[93] [9]), .C2(n_1_1_1155), .ZN(n_1_1_599));
   NAND3_X1 i_1_1_610 (.A1(n_1_1_603), .A2(n_1_1_602), .A3(n_1_1_601), .ZN(
      n_1_1_600));
   AOI22_X1 i_1_1_611 (.A1(\mem[11] [9]), .A2(n_1_1_1063), .B1(n_1_1_1035), 
      .B2(\mem[50] [9]), .ZN(n_1_1_601));
   AOI22_X1 i_1_1_612 (.A1(\mem[86] [9]), .A2(n_1_1_1142), .B1(n_1_1_1071), 
      .B2(\mem[5] [9]), .ZN(n_1_1_602));
   AOI22_X1 i_1_1_613 (.A1(\mem[54] [9]), .A2(n_1_1_1106), .B1(n_1_1_1025), 
      .B2(\mem[43] [9]), .ZN(n_1_1_603));
   AOI221_X1 i_1_1_614 (.A(n_1_1_605), .B1(n_1_1_1092), .B2(\mem[33] [9]), 
      .C1(\mem[91] [9]), .C2(n_1_1_1037), .ZN(n_1_1_604));
   NAND4_X1 i_1_1_615 (.A1(read_signal), .A2(n_1_1_608), .A3(n_1_1_607), 
      .A4(n_1_1_606), .ZN(n_1_1_605));
   AOI22_X1 i_1_1_616 (.A1(\mem[75] [9]), .A2(n_1_1_1061), .B1(n_1_1_1048), 
      .B2(\mem[10] [9]), .ZN(n_1_1_606));
   AOI22_X1 i_1_1_617 (.A1(\mem[12] [9]), .A2(n_1_1_1042), .B1(n_1_1_1033), 
      .B2(\mem[42] [9]), .ZN(n_1_1_607));
   NOR4_X1 i_1_1_618 (.A1(n_1_1_623), .A2(n_1_1_618), .A3(n_1_1_613), .A4(
      n_1_1_609), .ZN(n_1_1_608));
   NAND4_X1 i_1_1_619 (.A1(n_1_1_639), .A2(n_1_1_612), .A3(n_1_1_611), .A4(
      n_1_1_610), .ZN(n_1_1_609));
   AOI22_X1 i_1_1_620 (.A1(\mem[35] [9]), .A2(n_1_1_1094), .B1(n_1_1_1049), 
      .B2(\mem[17] [9]), .ZN(n_1_1_610));
   AOI22_X1 i_1_1_621 (.A1(\mem[4] [9]), .A2(n_1_1_1070), .B1(n_1_1_1052), 
      .B2(\mem[23] [9]), .ZN(n_1_1_611));
   AOI22_X1 i_1_1_622 (.A1(\mem[92] [9]), .A2(n_1_1_1153), .B1(n_1_1_1027), 
      .B2(\mem[27] [9]), .ZN(n_1_1_612));
   NAND4_X1 i_1_1_623 (.A1(n_1_1_617), .A2(n_1_1_616), .A3(n_1_1_615), .A4(
      n_1_1_614), .ZN(n_1_1_613));
   AOI22_X1 i_1_1_624 (.A1(\mem[97] [9]), .A2(n_1_1_1165), .B1(n_1_1_1026), 
      .B2(\mem[56] [9]), .ZN(n_1_1_614));
   AOI22_X1 i_1_1_625 (.A1(\mem[48] [9]), .A2(n_1_1_1104), .B1(n_1_1_1062), 
      .B2(\mem[84] [9]), .ZN(n_1_1_615));
   AOI22_X1 i_1_1_626 (.A1(\mem[77] [9]), .A2(n_1_1_1133), .B1(n_1_1_1038), 
      .B2(\mem[15] [9]), .ZN(n_1_1_616));
   AOI22_X1 i_1_1_627 (.A1(\mem[38] [9]), .A2(n_1_1_1097), .B1(n_1_1_1066), 
      .B2(\mem[0] [9]), .ZN(n_1_1_617));
   NAND4_X1 i_1_1_628 (.A1(n_1_1_622), .A2(n_1_1_621), .A3(n_1_1_620), .A4(
      n_1_1_619), .ZN(n_1_1_618));
   AOI22_X1 i_1_1_629 (.A1(\mem[47] [9]), .A2(n_1_1_1102), .B1(n_1_1_1032), 
      .B2(\mem[44] [9]), .ZN(n_1_1_619));
   AOI22_X1 i_1_1_630 (.A1(\mem[98] [9]), .A2(n_1_1_1168), .B1(n_1_1_1148), 
      .B2(\mem[89] [9]), .ZN(n_1_1_620));
   AOI22_X1 i_1_1_631 (.A1(\mem[65] [9]), .A2(n_1_1_1119), .B1(n_1_1_1029), 
      .B2(\mem[62] [9]), .ZN(n_1_1_621));
   AOI22_X1 i_1_1_632 (.A1(\mem[69] [9]), .A2(n_1_1_1123), .B1(n_1_1_1078), 
      .B2(\mem[16] [9]), .ZN(n_1_1_622));
   NAND4_X1 i_1_1_633 (.A1(n_1_1_627), .A2(n_1_1_626), .A3(n_1_1_625), .A4(
      n_1_1_624), .ZN(n_1_1_623));
   AOI22_X1 i_1_1_634 (.A1(\mem[57] [9]), .A2(n_1_1_1108), .B1(n_1_1_1053), 
      .B2(\mem[95] [9]), .ZN(n_1_1_624));
   AOI22_X1 i_1_1_635 (.A1(\mem[24] [9]), .A2(n_1_1_1083), .B1(n_1_1_1069), 
      .B2(\mem[3] [9]), .ZN(n_1_1_625));
   AOI22_X1 i_1_1_636 (.A1(\mem[71] [9]), .A2(n_1_1_1126), .B1(n_1_1_1091), 
      .B2(\mem[32] [9]), .ZN(n_1_1_626));
   AOI22_X1 i_1_1_637 (.A1(\mem[74] [9]), .A2(n_1_1_1055), .B1(n_1_1_1051), 
      .B2(\mem[29] [9]), .ZN(n_1_1_627));
   AOI221_X1 i_1_1_638 (.A(n_1_1_629), .B1(n_1_1_1060), .B2(\mem[28] [9]), 
      .C1(\mem[37] [9]), .C2(n_1_1_1096), .ZN(n_1_1_628));
   NAND3_X1 i_1_1_639 (.A1(n_1_1_640), .A2(n_1_1_631), .A3(n_1_1_630), .ZN(
      n_1_1_629));
   AOI22_X1 i_1_1_640 (.A1(\mem[51] [9]), .A2(n_1_1_1059), .B1(n_1_1_1041), 
      .B2(\mem[7] [9]), .ZN(n_1_1_630));
   AOI22_X1 i_1_1_641 (.A1(\mem[46] [9]), .A2(n_1_1_1101), .B1(n_1_1_1036), 
      .B2(\mem[14] [9]), .ZN(n_1_1_631));
   AOI221_X1 i_1_1_642 (.A(n_1_1_633), .B1(n_1_1_1064), .B2(\mem[18] [9]), 
      .C1(\mem[66] [9]), .C2(n_1_1_1120), .ZN(n_1_1_632));
   NAND3_X1 i_1_1_643 (.A1(n_1_1_636), .A2(n_1_1_635), .A3(n_1_1_634), .ZN(
      n_1_1_633));
   AOI22_X1 i_1_1_644 (.A1(\mem[45] [9]), .A2(n_1_1_1045), .B1(n_1_1_1039), 
      .B2(\mem[76] [9]), .ZN(n_1_1_634));
   AOI22_X1 i_1_1_645 (.A1(\mem[36] [9]), .A2(n_1_1_1095), .B1(n_1_1_1080), 
      .B2(\mem[19] [9]), .ZN(n_1_1_635));
   AOI22_X1 i_1_1_646 (.A1(\mem[40] [9]), .A2(n_1_1_1099), .B1(n_1_1_1058), 
      .B2(\mem[85] [9]), .ZN(n_1_1_636));
   AOI222_X1 i_1_1_647 (.A1(\mem[58] [9]), .A2(n_1_1_1109), .B1(n_1_1_1087), 
      .B2(\mem[30] [9]), .C1(n_1_1_1031), .C2(\mem[39] [9]), .ZN(n_1_1_637));
   AOI22_X1 i_1_1_648 (.A1(\mem[26] [9]), .A2(n_1_1_1044), .B1(n_1_1_1028), 
      .B2(\mem[82] [9]), .ZN(n_1_1_638));
   AOI22_X1 i_1_1_649 (.A1(\mem[67] [9]), .A2(n_1_1_1121), .B1(n_1_1_1050), 
      .B2(\mem[90] [9]), .ZN(n_1_1_639));
   AOI22_X1 i_1_1_650 (.A1(\mem[78] [9]), .A2(n_1_1_1134), .B1(n_1_1_1068), 
      .B2(\mem[2] [9]), .ZN(n_1_1_640));
   MUX2_X1 i_1_1_651 (.A(dataout[10]), .B(n_1_1_641), .S(read_signal), .Z(n_1_10));
   NAND4_X1 i_1_1_652 (.A1(n_1_1_684), .A2(n_1_1_679), .A3(n_1_1_660), .A4(
      n_1_1_642), .ZN(n_1_1_641));
   NOR4_X1 i_1_1_653 (.A1(n_1_1_655), .A2(n_1_1_651), .A3(n_1_1_646), .A4(
      n_1_1_643), .ZN(n_1_1_642));
   NAND4_X1 i_1_1_654 (.A1(n_1_1_703), .A2(n_1_1_699), .A3(n_1_1_645), .A4(
      n_1_1_644), .ZN(n_1_1_643));
   AOI22_X1 i_1_1_655 (.A1(\mem[70] [10]), .A2(n_1_1_1125), .B1(n_1_1_1057), 
      .B2(\mem[61] [10]), .ZN(n_1_1_644));
   AOI22_X1 i_1_1_656 (.A1(\mem[72] [10]), .A2(n_1_1_1127), .B1(n_1_1_1047), 
      .B2(\mem[83] [10]), .ZN(n_1_1_645));
   NAND4_X1 i_1_1_657 (.A1(n_1_1_650), .A2(n_1_1_649), .A3(n_1_1_648), .A4(
      n_1_1_647), .ZN(n_1_1_646));
   AOI22_X1 i_1_1_658 (.A1(\mem[73] [10]), .A2(n_1_1_1129), .B1(n_1_1_1062), 
      .B2(\mem[84] [10]), .ZN(n_1_1_647));
   AOI22_X1 i_1_1_659 (.A1(\mem[32] [10]), .A2(n_1_1_1091), .B1(n_1_1_1042), 
      .B2(\mem[12] [10]), .ZN(n_1_1_648));
   AOI22_X1 i_1_1_660 (.A1(\mem[100] [10]), .A2(n_1_1_1174), .B1(n_1_1_1126), 
      .B2(\mem[71] [10]), .ZN(n_1_1_649));
   AOI22_X1 i_1_1_661 (.A1(\mem[86] [10]), .A2(n_1_1_1142), .B1(n_1_1_1067), 
      .B2(\mem[1] [10]), .ZN(n_1_1_650));
   NAND4_X1 i_1_1_662 (.A1(n_1_1_700), .A2(n_1_1_654), .A3(n_1_1_653), .A4(
      n_1_1_652), .ZN(n_1_1_651));
   AOI22_X1 i_1_1_663 (.A1(\mem[38] [10]), .A2(n_1_1_1097), .B1(n_1_1_1060), 
      .B2(\mem[28] [10]), .ZN(n_1_1_652));
   AOI22_X1 i_1_1_664 (.A1(\mem[99] [10]), .A2(n_1_1_1171), .B1(n_1_1_1163), 
      .B2(\mem[96] [10]), .ZN(n_1_1_653));
   AOI22_X1 i_1_1_665 (.A1(\mem[19] [10]), .A2(n_1_1_1080), .B1(n_1_1_1078), 
      .B2(\mem[16] [10]), .ZN(n_1_1_654));
   NAND4_X1 i_1_1_666 (.A1(n_1_1_659), .A2(n_1_1_658), .A3(n_1_1_657), .A4(
      n_1_1_656), .ZN(n_1_1_655));
   AOI22_X1 i_1_1_667 (.A1(\mem[14] [10]), .A2(n_1_1_1036), .B1(n_1_1_1035), 
      .B2(\mem[50] [10]), .ZN(n_1_1_656));
   AOI22_X1 i_1_1_668 (.A1(\mem[46] [10]), .A2(n_1_1_1101), .B1(n_1_1_1043), 
      .B2(\mem[53] [10]), .ZN(n_1_1_657));
   AOI22_X1 i_1_1_669 (.A1(\mem[64] [10]), .A2(n_1_1_1118), .B1(n_1_1_1041), 
      .B2(\mem[7] [10]), .ZN(n_1_1_658));
   AOI22_X1 i_1_1_670 (.A1(\mem[63] [10]), .A2(n_1_1_1116), .B1(n_1_1_1048), 
      .B2(\mem[10] [10]), .ZN(n_1_1_659));
   NOR4_X1 i_1_1_671 (.A1(n_1_1_675), .A2(n_1_1_670), .A3(n_1_1_666), .A4(
      n_1_1_661), .ZN(n_1_1_660));
   NAND4_X1 i_1_1_672 (.A1(n_1_1_665), .A2(n_1_1_664), .A3(n_1_1_663), .A4(
      n_1_1_662), .ZN(n_1_1_661));
   AOI22_X1 i_1_1_673 (.A1(\mem[33] [10]), .A2(n_1_1_1092), .B1(n_1_1_1055), 
      .B2(\mem[74] [10]), .ZN(n_1_1_662));
   AOI22_X1 i_1_1_674 (.A1(\mem[47] [10]), .A2(n_1_1_1102), .B1(n_1_1_1083), 
      .B2(\mem[24] [10]), .ZN(n_1_1_663));
   AOI22_X1 i_1_1_675 (.A1(\mem[80] [10]), .A2(n_1_1_1138), .B1(n_1_1_1095), 
      .B2(\mem[36] [10]), .ZN(n_1_1_664));
   AOI22_X1 i_1_1_676 (.A1(\mem[90] [10]), .A2(n_1_1_1050), .B1(n_1_1_1044), 
      .B2(\mem[26] [10]), .ZN(n_1_1_665));
   NAND4_X1 i_1_1_677 (.A1(n_1_1_701), .A2(n_1_1_669), .A3(n_1_1_668), .A4(
      n_1_1_667), .ZN(n_1_1_666));
   AOI22_X1 i_1_1_678 (.A1(\mem[9] [10]), .A2(n_1_1_1074), .B1(n_1_1_1027), 
      .B2(\mem[27] [10]), .ZN(n_1_1_667));
   AOI22_X1 i_1_1_679 (.A1(\mem[66] [10]), .A2(n_1_1_1120), .B1(n_1_1_1073), 
      .B2(\mem[8] [10]), .ZN(n_1_1_668));
   AOI22_X1 i_1_1_680 (.A1(\mem[21] [10]), .A2(n_1_1_1081), .B1(n_1_1_1025), 
      .B2(\mem[43] [10]), .ZN(n_1_1_669));
   NAND4_X1 i_1_1_681 (.A1(n_1_1_674), .A2(n_1_1_673), .A3(n_1_1_672), .A4(
      n_1_1_671), .ZN(n_1_1_670));
   AOI22_X1 i_1_1_682 (.A1(\mem[97] [10]), .A2(n_1_1_1165), .B1(n_1_1_1104), 
      .B2(\mem[48] [10]), .ZN(n_1_1_671));
   AOI22_X1 i_1_1_683 (.A1(\mem[69] [10]), .A2(n_1_1_1123), .B1(n_1_1_1063), 
      .B2(\mem[11] [10]), .ZN(n_1_1_672));
   AOI22_X1 i_1_1_684 (.A1(\mem[94] [10]), .A2(n_1_1_1157), .B1(n_1_1_1053), 
      .B2(\mem[95] [10]), .ZN(n_1_1_673));
   AOI22_X1 i_1_1_685 (.A1(\mem[2] [10]), .A2(n_1_1_1068), .B1(n_1_1_1038), 
      .B2(\mem[15] [10]), .ZN(n_1_1_674));
   NAND4_X1 i_1_1_686 (.A1(n_1_1_704), .A2(n_1_1_678), .A3(n_1_1_677), .A4(
      n_1_1_676), .ZN(n_1_1_675));
   AOI22_X1 i_1_1_687 (.A1(\mem[92] [10]), .A2(n_1_1_1153), .B1(n_1_1_1087), 
      .B2(\mem[30] [10]), .ZN(n_1_1_676));
   AOI22_X1 i_1_1_688 (.A1(\mem[89] [10]), .A2(n_1_1_1148), .B1(n_1_1_1051), 
      .B2(\mem[29] [10]), .ZN(n_1_1_677));
   AOI22_X1 i_1_1_689 (.A1(\mem[57] [10]), .A2(n_1_1_1108), .B1(n_1_1_1106), 
      .B2(\mem[54] [10]), .ZN(n_1_1_678));
   AOI221_X1 i_1_1_690 (.A(n_1_1_680), .B1(n_1_1_1109), .B2(\mem[58] [10]), 
      .C1(\mem[82] [10]), .C2(n_1_1_1028), .ZN(n_1_1_679));
   NAND4_X1 i_1_1_691 (.A1(n_1_1_705), .A2(n_1_1_683), .A3(n_1_1_682), .A4(
      n_1_1_681), .ZN(n_1_1_680));
   AOI22_X1 i_1_1_692 (.A1(\mem[41] [10]), .A2(n_1_1_1100), .B1(n_1_1_1075), 
      .B2(\mem[13] [10]), .ZN(n_1_1_681));
   AOI22_X1 i_1_1_693 (.A1(\mem[68] [10]), .A2(n_1_1_1122), .B1(n_1_1_1033), 
      .B2(\mem[42] [10]), .ZN(n_1_1_682));
   AOI22_X1 i_1_1_694 (.A1(\mem[44] [10]), .A2(n_1_1_1032), .B1(n_1_1_1030), 
      .B2(\mem[20] [10]), .ZN(n_1_1_683));
   AOI221_X1 i_1_1_695 (.A(n_1_1_685), .B1(n_1_1_1093), .B2(\mem[34] [10]), 
      .C1(\mem[65] [10]), .C2(n_1_1_1119), .ZN(n_1_1_684));
   NAND4_X1 i_1_1_696 (.A1(n_1_1_698), .A2(n_1_1_693), .A3(n_1_1_687), .A4(
      n_1_1_686), .ZN(n_1_1_685));
   AOI22_X1 i_1_1_697 (.A1(\mem[91] [10]), .A2(n_1_1_1037), .B1(n_1_1_1026), 
      .B2(\mem[56] [10]), .ZN(n_1_1_686));
   AOI221_X1 i_1_1_698 (.A(n_1_1_688), .B1(n_1_1_1072), .B2(\mem[6] [10]), 
      .C1(\mem[60] [10]), .C2(n_1_1_1046), .ZN(n_1_1_687));
   NAND4_X1 i_1_1_699 (.A1(n_1_1_692), .A2(n_1_1_691), .A3(n_1_1_690), .A4(
      n_1_1_689), .ZN(n_1_1_688));
   AOI22_X1 i_1_1_700 (.A1(\mem[98] [10]), .A2(n_1_1_1168), .B1(n_1_1_1071), 
      .B2(\mem[5] [10]), .ZN(n_1_1_689));
   AOI22_X1 i_1_1_701 (.A1(\mem[35] [10]), .A2(n_1_1_1094), .B1(n_1_1_1061), 
      .B2(\mem[75] [10]), .ZN(n_1_1_690));
   AOI22_X1 i_1_1_702 (.A1(\mem[77] [10]), .A2(n_1_1_1133), .B1(n_1_1_1056), 
      .B2(\mem[88] [10]), .ZN(n_1_1_691));
   AOI22_X1 i_1_1_703 (.A1(\mem[25] [10]), .A2(n_1_1_1084), .B1(n_1_1_1054), 
      .B2(\mem[22] [10]), .ZN(n_1_1_692));
   AOI221_X1 i_1_1_704 (.A(n_1_1_694), .B1(n_1_1_1052), .B2(\mem[23] [10]), 
      .C1(\mem[79] [10]), .C2(n_1_1_1135), .ZN(n_1_1_693));
   NAND4_X1 i_1_1_705 (.A1(n_1_1_702), .A2(n_1_1_697), .A3(n_1_1_696), .A4(
      n_1_1_695), .ZN(n_1_1_694));
   AOI22_X1 i_1_1_706 (.A1(\mem[59] [10]), .A2(n_1_1_1111), .B1(n_1_1_1040), 
      .B2(\mem[52] [10]), .ZN(n_1_1_695));
   AOI22_X1 i_1_1_707 (.A1(\mem[87] [10]), .A2(n_1_1_1144), .B1(n_1_1_1070), 
      .B2(\mem[4] [10]), .ZN(n_1_1_696));
   AOI22_X1 i_1_1_708 (.A1(\mem[78] [10]), .A2(n_1_1_1134), .B1(n_1_1_1069), 
      .B2(\mem[3] [10]), .ZN(n_1_1_697));
   AOI222_X1 i_1_1_709 (.A1(\mem[67] [10]), .A2(n_1_1_1121), .B1(n_1_1_1096), 
      .B2(\mem[37] [10]), .C1(n_1_1_1059), .C2(\mem[51] [10]), .ZN(n_1_1_698));
   AOI22_X1 i_1_1_710 (.A1(\mem[49] [10]), .A2(n_1_1_1105), .B1(n_1_1_1066), 
      .B2(\mem[0] [10]), .ZN(n_1_1_699));
   AOI22_X1 i_1_1_711 (.A1(\mem[18] [10]), .A2(n_1_1_1064), .B1(n_1_1_1045), 
      .B2(\mem[45] [10]), .ZN(n_1_1_700));
   AOI22_X1 i_1_1_712 (.A1(\mem[85] [10]), .A2(n_1_1_1058), .B1(n_1_1_1029), 
      .B2(\mem[62] [10]), .ZN(n_1_1_701));
   AOI22_X1 i_1_1_713 (.A1(\mem[81] [10]), .A2(n_1_1_1139), .B1(n_1_1_1031), 
      .B2(\mem[39] [10]), .ZN(n_1_1_702));
   AOI22_X1 i_1_1_714 (.A1(\mem[93] [10]), .A2(n_1_1_1155), .B1(n_1_1_1099), 
      .B2(\mem[40] [10]), .ZN(n_1_1_703));
   AOI22_X1 i_1_1_715 (.A1(\mem[17] [10]), .A2(n_1_1_1049), .B1(n_1_1_1039), 
      .B2(\mem[76] [10]), .ZN(n_1_1_704));
   AOI22_X1 i_1_1_716 (.A1(\mem[55] [10]), .A2(n_1_1_1107), .B1(n_1_1_1088), 
      .B2(\mem[31] [10]), .ZN(n_1_1_705));
   MUX2_X1 i_1_1_717 (.A(dataout[11]), .B(n_1_1_706), .S(read_signal), .Z(n_1_11));
   NAND4_X1 i_1_1_718 (.A1(n_1_1_722), .A2(n_1_1_717), .A3(n_1_1_712), .A4(
      n_1_1_707), .ZN(n_1_1_706));
   AOI221_X1 i_1_1_719 (.A(n_1_1_708), .B1(n_1_1_1049), .B2(\mem[17] [11]), 
      .C1(\mem[97] [11]), .C2(n_1_1_1165), .ZN(n_1_1_707));
   NAND3_X1 i_1_1_720 (.A1(n_1_1_711), .A2(n_1_1_710), .A3(n_1_1_709), .ZN(
      n_1_1_708));
   AOI22_X1 i_1_1_721 (.A1(\mem[64] [11]), .A2(n_1_1_1118), .B1(n_1_1_1069), 
      .B2(\mem[3] [11]), .ZN(n_1_1_709));
   AOI22_X1 i_1_1_722 (.A1(\mem[10] [11]), .A2(n_1_1_1048), .B1(n_1_1_1038), 
      .B2(\mem[15] [11]), .ZN(n_1_1_710));
   AOI22_X1 i_1_1_723 (.A1(\mem[92] [11]), .A2(n_1_1_1153), .B1(n_1_1_1063), 
      .B2(\mem[11] [11]), .ZN(n_1_1_711));
   AOI221_X1 i_1_1_724 (.A(n_1_1_713), .B1(n_1_1_1032), .B2(\mem[44] [11]), 
      .C1(\mem[52] [11]), .C2(n_1_1_1040), .ZN(n_1_1_712));
   NAND3_X1 i_1_1_725 (.A1(n_1_1_716), .A2(n_1_1_715), .A3(n_1_1_714), .ZN(
      n_1_1_713));
   AOI22_X1 i_1_1_726 (.A1(\mem[46] [11]), .A2(n_1_1_1101), .B1(n_1_1_1036), 
      .B2(\mem[14] [11]), .ZN(n_1_1_714));
   AOI22_X1 i_1_1_727 (.A1(\mem[63] [11]), .A2(n_1_1_1116), .B1(n_1_1_1026), 
      .B2(\mem[56] [11]), .ZN(n_1_1_715));
   AOI22_X1 i_1_1_728 (.A1(\mem[57] [11]), .A2(n_1_1_1108), .B1(n_1_1_1096), 
      .B2(\mem[37] [11]), .ZN(n_1_1_716));
   AOI221_X1 i_1_1_729 (.A(n_1_1_718), .B1(n_1_1_1133), .B2(\mem[77] [11]), 
      .C1(\mem[85] [11]), .C2(n_1_1_1058), .ZN(n_1_1_717));
   NAND3_X1 i_1_1_730 (.A1(n_1_1_721), .A2(n_1_1_720), .A3(n_1_1_719), .ZN(
      n_1_1_718));
   AOI22_X1 i_1_1_731 (.A1(\mem[87] [11]), .A2(n_1_1_1144), .B1(n_1_1_1064), 
      .B2(\mem[18] [11]), .ZN(n_1_1_719));
   AOI22_X1 i_1_1_732 (.A1(\mem[55] [11]), .A2(n_1_1_1107), .B1(n_1_1_1043), 
      .B2(\mem[53] [11]), .ZN(n_1_1_720));
   AOI22_X1 i_1_1_733 (.A1(\mem[68] [11]), .A2(n_1_1_1122), .B1(n_1_1_1052), 
      .B2(\mem[23] [11]), .ZN(n_1_1_721));
   NOR4_X1 i_1_1_734 (.A1(n_1_1_738), .A2(n_1_1_737), .A3(n_1_1_731), .A4(
      n_1_1_723), .ZN(n_1_1_722));
   NAND3_X1 i_1_1_735 (.A1(n_1_1_755), .A2(n_1_1_730), .A3(n_1_1_724), .ZN(
      n_1_1_723));
   AOI221_X1 i_1_1_736 (.A(n_1_1_725), .B1(n_1_1_1105), .B2(\mem[49] [11]), 
      .C1(\mem[78] [11]), .C2(n_1_1_1134), .ZN(n_1_1_724));
   NAND4_X1 i_1_1_737 (.A1(n_1_1_729), .A2(n_1_1_728), .A3(n_1_1_727), .A4(
      n_1_1_726), .ZN(n_1_1_725));
   AOI22_X1 i_1_1_738 (.A1(\mem[19] [11]), .A2(n_1_1_1080), .B1(n_1_1_1072), 
      .B2(\mem[6] [11]), .ZN(n_1_1_726));
   AOI22_X1 i_1_1_739 (.A1(\mem[5] [11]), .A2(n_1_1_1071), .B1(n_1_1_1061), 
      .B2(\mem[75] [11]), .ZN(n_1_1_727));
   AOI22_X1 i_1_1_740 (.A1(\mem[99] [11]), .A2(n_1_1_1171), .B1(n_1_1_1084), 
      .B2(\mem[25] [11]), .ZN(n_1_1_728));
   AOI22_X1 i_1_1_741 (.A1(\mem[84] [11]), .A2(n_1_1_1062), .B1(n_1_1_1041), 
      .B2(\mem[7] [11]), .ZN(n_1_1_729));
   AOI222_X1 i_1_1_742 (.A1(\mem[59] [11]), .A2(n_1_1_1111), .B1(n_1_1_1074), 
      .B2(\mem[9] [11]), .C1(n_1_1_1066), .C2(\mem[0] [11]), .ZN(n_1_1_730));
   NAND4_X1 i_1_1_743 (.A1(n_1_1_735), .A2(n_1_1_734), .A3(n_1_1_733), .A4(
      n_1_1_732), .ZN(n_1_1_731));
   AOI222_X1 i_1_1_744 (.A1(\mem[89] [11]), .A2(n_1_1_1148), .B1(n_1_1_1125), 
      .B2(\mem[70] [11]), .C1(n_1_1_1028), .C2(\mem[82] [11]), .ZN(n_1_1_732));
   AOI22_X1 i_1_1_745 (.A1(\mem[81] [11]), .A2(n_1_1_1139), .B1(n_1_1_1093), 
      .B2(\mem[34] [11]), .ZN(n_1_1_733));
   AOI222_X1 i_1_1_746 (.A1(\mem[98] [11]), .A2(n_1_1_1168), .B1(n_1_1_1155), 
      .B2(\mem[93] [11]), .C1(n_1_1_1054), .C2(\mem[22] [11]), .ZN(n_1_1_734));
   AOI221_X1 i_1_1_747 (.A(n_1_1_736), .B1(n_1_1_1060), .B2(\mem[28] [11]), 
      .C1(\mem[73] [11]), .C2(n_1_1_1129), .ZN(n_1_1_735));
   NAND3_X1 i_1_1_748 (.A1(n_1_1_767), .A2(n_1_1_763), .A3(n_1_1_751), .ZN(
      n_1_1_736));
   NAND4_X1 i_1_1_749 (.A1(n_1_1_760), .A2(n_1_1_759), .A3(n_1_1_750), .A4(
      n_1_1_749), .ZN(n_1_1_737));
   NAND4_X1 i_1_1_750 (.A1(n_1_1_766), .A2(n_1_1_754), .A3(n_1_1_746), .A4(
      n_1_1_739), .ZN(n_1_1_738));
   NOR4_X1 i_1_1_751 (.A1(n_1_1_743), .A2(n_1_1_742), .A3(n_1_1_741), .A4(
      n_1_1_740), .ZN(n_1_1_739));
   NAND4_X1 i_1_1_752 (.A1(n_1_1_769), .A2(n_1_1_764), .A3(n_1_1_758), .A4(
      n_1_1_745), .ZN(n_1_1_740));
   NAND4_X1 i_1_1_753 (.A1(n_1_1_770), .A2(n_1_1_768), .A3(n_1_1_748), .A4(
      n_1_1_747), .ZN(n_1_1_741));
   NAND4_X1 i_1_1_754 (.A1(n_1_1_765), .A2(n_1_1_761), .A3(n_1_1_753), .A4(
      n_1_1_752), .ZN(n_1_1_742));
   NAND4_X1 i_1_1_755 (.A1(n_1_1_762), .A2(n_1_1_757), .A3(n_1_1_756), .A4(
      n_1_1_744), .ZN(n_1_1_743));
   AOI22_X1 i_1_1_756 (.A1(\mem[36] [11]), .A2(n_1_1_1095), .B1(n_1_1_1037), 
      .B2(\mem[91] [11]), .ZN(n_1_1_744));
   AOI22_X1 i_1_1_757 (.A1(\mem[65] [11]), .A2(n_1_1_1119), .B1(n_1_1_1029), 
      .B2(\mem[62] [11]), .ZN(n_1_1_745));
   AOI22_X1 i_1_1_758 (.A1(\mem[30] [11]), .A2(n_1_1_1087), .B1(n_1_1_1056), 
      .B2(\mem[88] [11]), .ZN(n_1_1_746));
   AOI22_X1 i_1_1_759 (.A1(\mem[66] [11]), .A2(n_1_1_1120), .B1(n_1_1_1100), 
      .B2(\mem[41] [11]), .ZN(n_1_1_747));
   AOI22_X1 i_1_1_760 (.A1(\mem[94] [11]), .A2(n_1_1_1157), .B1(n_1_1_1078), 
      .B2(\mem[16] [11]), .ZN(n_1_1_748));
   AOI22_X1 i_1_1_761 (.A1(\mem[45] [11]), .A2(n_1_1_1045), .B1(n_1_1_1031), 
      .B2(\mem[39] [11]), .ZN(n_1_1_749));
   AOI22_X1 i_1_1_762 (.A1(\mem[31] [11]), .A2(n_1_1_1088), .B1(n_1_1_1030), 
      .B2(\mem[20] [11]), .ZN(n_1_1_750));
   AOI22_X1 i_1_1_763 (.A1(\mem[79] [11]), .A2(n_1_1_1135), .B1(n_1_1_1042), 
      .B2(\mem[12] [11]), .ZN(n_1_1_751));
   AOI22_X1 i_1_1_764 (.A1(\mem[69] [11]), .A2(n_1_1_1123), .B1(n_1_1_1104), 
      .B2(\mem[48] [11]), .ZN(n_1_1_752));
   AOI22_X1 i_1_1_765 (.A1(\mem[72] [11]), .A2(n_1_1_1127), .B1(n_1_1_1073), 
      .B2(\mem[8] [11]), .ZN(n_1_1_753));
   AOI22_X1 i_1_1_766 (.A1(\mem[35] [11]), .A2(n_1_1_1094), .B1(n_1_1_1091), 
      .B2(\mem[32] [11]), .ZN(n_1_1_754));
   AOI22_X1 i_1_1_767 (.A1(\mem[51] [11]), .A2(n_1_1_1059), .B1(n_1_1_1025), 
      .B2(\mem[43] [11]), .ZN(n_1_1_755));
   AOI22_X1 i_1_1_768 (.A1(\mem[38] [11]), .A2(n_1_1_1097), .B1(n_1_1_1053), 
      .B2(\mem[95] [11]), .ZN(n_1_1_756));
   AOI22_X1 i_1_1_769 (.A1(\mem[74] [11]), .A2(n_1_1_1055), .B1(n_1_1_1044), 
      .B2(\mem[26] [11]), .ZN(n_1_1_757));
   AOI22_X1 i_1_1_770 (.A1(\mem[1] [11]), .A2(n_1_1_1067), .B1(n_1_1_1057), 
      .B2(\mem[61] [11]), .ZN(n_1_1_758));
   AOI22_X1 i_1_1_771 (.A1(\mem[71] [11]), .A2(n_1_1_1126), .B1(n_1_1_1102), 
      .B2(\mem[47] [11]), .ZN(n_1_1_759));
   AOI22_X1 i_1_1_772 (.A1(\mem[96] [11]), .A2(n_1_1_1163), .B1(n_1_1_1070), 
      .B2(\mem[4] [11]), .ZN(n_1_1_760));
   AOI22_X1 i_1_1_773 (.A1(\mem[21] [11]), .A2(n_1_1_1081), .B1(n_1_1_1027), 
      .B2(\mem[27] [11]), .ZN(n_1_1_761));
   AOI22_X1 i_1_1_774 (.A1(\mem[80] [11]), .A2(n_1_1_1138), .B1(n_1_1_1106), 
      .B2(\mem[54] [11]), .ZN(n_1_1_762));
   AOI22_X1 i_1_1_775 (.A1(\mem[100] [11]), .A2(n_1_1_1174), .B1(n_1_1_1051), 
      .B2(\mem[29] [11]), .ZN(n_1_1_763));
   AOI22_X1 i_1_1_776 (.A1(\mem[76] [11]), .A2(n_1_1_1039), .B1(n_1_1_1035), 
      .B2(\mem[50] [11]), .ZN(n_1_1_764));
   AOI22_X1 i_1_1_777 (.A1(\mem[58] [11]), .A2(n_1_1_1109), .B1(n_1_1_1083), 
      .B2(\mem[24] [11]), .ZN(n_1_1_765));
   AOI22_X1 i_1_1_778 (.A1(\mem[40] [11]), .A2(n_1_1_1099), .B1(n_1_1_1046), 
      .B2(\mem[60] [11]), .ZN(n_1_1_766));
   AOI22_X1 i_1_1_779 (.A1(\mem[2] [11]), .A2(n_1_1_1068), .B1(n_1_1_1047), 
      .B2(\mem[83] [11]), .ZN(n_1_1_767));
   AOI22_X1 i_1_1_780 (.A1(\mem[90] [11]), .A2(n_1_1_1050), .B1(n_1_1_1033), 
      .B2(\mem[42] [11]), .ZN(n_1_1_768));
   AOI22_X1 i_1_1_781 (.A1(\mem[86] [11]), .A2(n_1_1_1142), .B1(n_1_1_1121), 
      .B2(\mem[67] [11]), .ZN(n_1_1_769));
   AOI22_X1 i_1_1_782 (.A1(\mem[33] [11]), .A2(n_1_1_1092), .B1(n_1_1_1075), 
      .B2(\mem[13] [11]), .ZN(n_1_1_770));
   MUX2_X1 i_1_1_783 (.A(dataout[12]), .B(n_1_1_771), .S(read_signal), .Z(n_1_12));
   NAND4_X1 i_1_1_784 (.A1(n_1_1_795), .A2(n_1_1_774), .A3(n_1_1_773), .A4(
      n_1_1_772), .ZN(n_1_1_771));
   AOI222_X1 i_1_1_785 (.A1(\mem[96] [12]), .A2(n_1_1_1163), .B1(n_1_1_1100), 
      .B2(\mem[41] [12]), .C1(n_1_1_1088), .C2(\mem[31] [12]), .ZN(n_1_1_772));
   AOI22_X1 i_1_1_786 (.A1(\mem[37] [12]), .A2(n_1_1_1096), .B1(n_1_1_1032), 
      .B2(\mem[44] [12]), .ZN(n_1_1_773));
   NOR4_X1 i_1_1_787 (.A1(n_1_1_788), .A2(n_1_1_779), .A3(n_1_1_778), .A4(
      n_1_1_775), .ZN(n_1_1_774));
   NAND4_X1 i_1_1_788 (.A1(n_1_1_826), .A2(n_1_1_818), .A3(n_1_1_777), .A4(
      n_1_1_776), .ZN(n_1_1_775));
   AOI22_X1 i_1_1_789 (.A1(\mem[71] [12]), .A2(n_1_1_1126), .B1(n_1_1_1080), 
      .B2(\mem[19] [12]), .ZN(n_1_1_776));
   AOI22_X1 i_1_1_790 (.A1(\mem[69] [12]), .A2(n_1_1_1123), .B1(n_1_1_1097), 
      .B2(\mem[38] [12]), .ZN(n_1_1_777));
   NAND4_X1 i_1_1_791 (.A1(n_1_1_825), .A2(n_1_1_822), .A3(n_1_1_821), .A4(
      n_1_1_816), .ZN(n_1_1_778));
   NAND4_X1 i_1_1_792 (.A1(n_1_1_787), .A2(n_1_1_783), .A3(n_1_1_782), .A4(
      n_1_1_780), .ZN(n_1_1_779));
   AOI221_X1 i_1_1_793 (.A(n_1_1_781), .B1(n_1_1_1094), .B2(\mem[35] [12]), 
      .C1(\mem[63] [12]), .C2(n_1_1_1116), .ZN(n_1_1_780));
   NAND4_X1 i_1_1_794 (.A1(n_1_1_832), .A2(n_1_1_824), .A3(n_1_1_823), .A4(
      n_1_1_817), .ZN(n_1_1_781));
   AOI222_X1 i_1_1_795 (.A1(\mem[64] [12]), .A2(n_1_1_1118), .B1(n_1_1_1043), 
      .B2(\mem[53] [12]), .C1(n_1_1_1026), .C2(\mem[56] [12]), .ZN(n_1_1_782));
   AOI21_X1 i_1_1_796 (.A(n_1_1_784), .B1(n_1_1_1040), .B2(\mem[52] [12]), 
      .ZN(n_1_1_783));
   NAND3_X1 i_1_1_797 (.A1(n_1_1_831), .A2(n_1_1_786), .A3(n_1_1_785), .ZN(
      n_1_1_784));
   AOI222_X1 i_1_1_798 (.A1(\mem[99] [12]), .A2(n_1_1_1171), .B1(n_1_1_1144), 
      .B2(\mem[87] [12]), .C1(n_1_1_1056), .C2(\mem[88] [12]), .ZN(n_1_1_785));
   AOI22_X1 i_1_1_799 (.A1(\mem[40] [12]), .A2(n_1_1_1099), .B1(n_1_1_1050), 
      .B2(\mem[90] [12]), .ZN(n_1_1_786));
   AOI22_X1 i_1_1_800 (.A1(\mem[68] [12]), .A2(n_1_1_1122), .B1(n_1_1_1038), 
      .B2(\mem[15] [12]), .ZN(n_1_1_787));
   NAND4_X1 i_1_1_801 (.A1(n_1_1_828), .A2(n_1_1_794), .A3(n_1_1_793), .A4(
      n_1_1_789), .ZN(n_1_1_788));
   AOI221_X1 i_1_1_802 (.A(n_1_1_790), .B1(n_1_1_1129), .B2(\mem[73] [12]), 
      .C1(\mem[95] [12]), .C2(n_1_1_1053), .ZN(n_1_1_789));
   NAND3_X1 i_1_1_803 (.A1(n_1_1_830), .A2(n_1_1_792), .A3(n_1_1_791), .ZN(
      n_1_1_790));
   AOI22_X1 i_1_1_804 (.A1(\mem[81] [12]), .A2(n_1_1_1139), .B1(n_1_1_1039), 
      .B2(\mem[76] [12]), .ZN(n_1_1_791));
   AOI22_X1 i_1_1_805 (.A1(\mem[57] [12]), .A2(n_1_1_1108), .B1(n_1_1_1048), 
      .B2(\mem[10] [12]), .ZN(n_1_1_792));
   AOI222_X1 i_1_1_806 (.A1(\mem[72] [12]), .A2(n_1_1_1127), .B1(n_1_1_1125), 
      .B2(\mem[70] [12]), .C1(n_1_1_1058), .C2(\mem[85] [12]), .ZN(n_1_1_793));
   AOI222_X1 i_1_1_807 (.A1(\mem[97] [12]), .A2(n_1_1_1165), .B1(n_1_1_1138), 
      .B2(\mem[80] [12]), .C1(n_1_1_1072), .C2(\mem[6] [12]), .ZN(n_1_1_794));
   AOI221_X1 i_1_1_808 (.A(n_1_1_796), .B1(n_1_1_1030), .B2(\mem[20] [12]), 
      .C1(\mem[93] [12]), .C2(n_1_1_1155), .ZN(n_1_1_795));
   NAND4_X1 i_1_1_809 (.A1(n_1_1_820), .A2(n_1_1_819), .A3(n_1_1_814), .A4(
      n_1_1_797), .ZN(n_1_1_796));
   NOR4_X1 i_1_1_810 (.A1(n_1_1_810), .A2(n_1_1_805), .A3(n_1_1_802), .A4(
      n_1_1_798), .ZN(n_1_1_797));
   NAND4_X1 i_1_1_811 (.A1(n_1_1_829), .A2(n_1_1_801), .A3(n_1_1_800), .A4(
      n_1_1_799), .ZN(n_1_1_798));
   AOI22_X1 i_1_1_812 (.A1(\mem[16] [12]), .A2(n_1_1_1078), .B1(n_1_1_1061), 
      .B2(\mem[75] [12]), .ZN(n_1_1_799));
   AOI22_X1 i_1_1_813 (.A1(\mem[92] [12]), .A2(n_1_1_1153), .B1(n_1_1_1107), 
      .B2(\mem[55] [12]), .ZN(n_1_1_800));
   AOI22_X1 i_1_1_814 (.A1(\mem[58] [12]), .A2(n_1_1_1109), .B1(n_1_1_1092), 
      .B2(\mem[33] [12]), .ZN(n_1_1_801));
   NAND3_X1 i_1_1_815 (.A1(n_1_1_815), .A2(n_1_1_804), .A3(n_1_1_803), .ZN(
      n_1_1_802));
   AOI222_X1 i_1_1_816 (.A1(\mem[54] [12]), .A2(n_1_1_1106), .B1(n_1_1_1093), 
      .B2(\mem[34] [12]), .C1(n_1_1_1075), .C2(\mem[13] [12]), .ZN(n_1_1_803));
   AOI222_X1 i_1_1_817 (.A1(\mem[25] [12]), .A2(n_1_1_1084), .B1(n_1_1_1036), 
      .B2(\mem[14] [12]), .C1(n_1_1_1033), .C2(\mem[42] [12]), .ZN(n_1_1_804));
   NAND4_X1 i_1_1_818 (.A1(n_1_1_809), .A2(n_1_1_808), .A3(n_1_1_807), .A4(
      n_1_1_806), .ZN(n_1_1_805));
   AOI22_X1 i_1_1_819 (.A1(\mem[21] [12]), .A2(n_1_1_1081), .B1(n_1_1_1068), 
      .B2(\mem[2] [12]), .ZN(n_1_1_806));
   AOI22_X1 i_1_1_820 (.A1(\mem[65] [12]), .A2(n_1_1_1119), .B1(n_1_1_1029), 
      .B2(\mem[62] [12]), .ZN(n_1_1_807));
   AOI22_X1 i_1_1_821 (.A1(\mem[98] [12]), .A2(n_1_1_1168), .B1(n_1_1_1071), 
      .B2(\mem[5] [12]), .ZN(n_1_1_808));
   AOI22_X1 i_1_1_822 (.A1(\mem[77] [12]), .A2(n_1_1_1133), .B1(n_1_1_1104), 
      .B2(\mem[48] [12]), .ZN(n_1_1_809));
   NAND4_X1 i_1_1_823 (.A1(n_1_1_827), .A2(n_1_1_813), .A3(n_1_1_812), .A4(
      n_1_1_811), .ZN(n_1_1_810));
   AOI22_X1 i_1_1_824 (.A1(\mem[30] [12]), .A2(n_1_1_1087), .B1(n_1_1_1055), 
      .B2(\mem[74] [12]), .ZN(n_1_1_811));
   AOI22_X1 i_1_1_825 (.A1(\mem[12] [12]), .A2(n_1_1_1042), .B1(n_1_1_1037), 
      .B2(\mem[91] [12]), .ZN(n_1_1_812));
   AOI22_X1 i_1_1_826 (.A1(\mem[100] [12]), .A2(n_1_1_1174), .B1(n_1_1_1051), 
      .B2(\mem[29] [12]), .ZN(n_1_1_813));
   AOI22_X1 i_1_1_827 (.A1(\mem[36] [12]), .A2(n_1_1_1095), .B1(n_1_1_1064), 
      .B2(\mem[18] [12]), .ZN(n_1_1_814));
   AOI22_X1 i_1_1_828 (.A1(\mem[1] [12]), .A2(n_1_1_1067), .B1(n_1_1_1062), 
      .B2(\mem[84] [12]), .ZN(n_1_1_815));
   AOI22_X1 i_1_1_829 (.A1(\mem[94] [12]), .A2(n_1_1_1157), .B1(n_1_1_1148), 
      .B2(\mem[89] [12]), .ZN(n_1_1_816));
   AOI22_X1 i_1_1_830 (.A1(\mem[79] [12]), .A2(n_1_1_1135), .B1(n_1_1_1073), 
      .B2(\mem[8] [12]), .ZN(n_1_1_817));
   AOI22_X1 i_1_1_831 (.A1(\mem[46] [12]), .A2(n_1_1_1101), .B1(n_1_1_1069), 
      .B2(\mem[3] [12]), .ZN(n_1_1_818));
   AOI22_X1 i_1_1_832 (.A1(\mem[17] [12]), .A2(n_1_1_1049), .B1(n_1_1_1035), 
      .B2(\mem[50] [12]), .ZN(n_1_1_819));
   AOI222_X1 i_1_1_833 (.A1(\mem[59] [12]), .A2(n_1_1_1111), .B1(n_1_1_1074), 
      .B2(\mem[9] [12]), .C1(n_1_1_1046), .C2(\mem[60] [12]), .ZN(n_1_1_820));
   AOI22_X1 i_1_1_834 (.A1(\mem[47] [12]), .A2(n_1_1_1102), .B1(n_1_1_1045), 
      .B2(\mem[45] [12]), .ZN(n_1_1_821));
   AOI22_X1 i_1_1_835 (.A1(\mem[66] [12]), .A2(n_1_1_1120), .B1(n_1_1_1059), 
      .B2(\mem[51] [12]), .ZN(n_1_1_822));
   AOI22_X1 i_1_1_836 (.A1(\mem[22] [12]), .A2(n_1_1_1054), .B1(n_1_1_1027), 
      .B2(\mem[27] [12]), .ZN(n_1_1_823));
   AOI22_X1 i_1_1_837 (.A1(\mem[49] [12]), .A2(n_1_1_1105), .B1(n_1_1_1063), 
      .B2(\mem[11] [12]), .ZN(n_1_1_824));
   AOI22_X1 i_1_1_838 (.A1(\mem[78] [12]), .A2(n_1_1_1134), .B1(n_1_1_1057), 
      .B2(\mem[61] [12]), .ZN(n_1_1_825));
   AOI22_X1 i_1_1_839 (.A1(\mem[7] [12]), .A2(n_1_1_1041), .B1(n_1_1_1025), 
      .B2(\mem[43] [12]), .ZN(n_1_1_826));
   AOI22_X1 i_1_1_840 (.A1(\mem[86] [12]), .A2(n_1_1_1142), .B1(n_1_1_1044), 
      .B2(\mem[26] [12]), .ZN(n_1_1_827));
   AOI22_X1 i_1_1_841 (.A1(\mem[32] [12]), .A2(n_1_1_1091), .B1(n_1_1_1066), 
      .B2(\mem[0] [12]), .ZN(n_1_1_828));
   AOI22_X1 i_1_1_842 (.A1(\mem[67] [12]), .A2(n_1_1_1121), .B1(n_1_1_1047), 
      .B2(\mem[83] [12]), .ZN(n_1_1_829));
   AOI22_X1 i_1_1_843 (.A1(\mem[24] [12]), .A2(n_1_1_1083), .B1(n_1_1_1060), 
      .B2(\mem[28] [12]), .ZN(n_1_1_830));
   AOI22_X1 i_1_1_844 (.A1(\mem[23] [12]), .A2(n_1_1_1052), .B1(n_1_1_1028), 
      .B2(\mem[82] [12]), .ZN(n_1_1_831));
   AOI22_X1 i_1_1_845 (.A1(\mem[4] [12]), .A2(n_1_1_1070), .B1(n_1_1_1031), 
      .B2(\mem[39] [12]), .ZN(n_1_1_832));
   MUX2_X1 i_1_1_846 (.A(dataout[13]), .B(n_1_1_833), .S(read_signal), .Z(n_1_13));
   NAND3_X1 i_1_1_847 (.A1(n_1_1_877), .A2(n_1_1_855), .A3(n_1_1_834), .ZN(
      n_1_1_833));
   NOR3_X1 i_1_1_848 (.A1(n_1_1_850), .A2(n_1_1_838), .A3(n_1_1_835), .ZN(
      n_1_1_834));
   NAND4_X1 i_1_1_849 (.A1(n_1_1_896), .A2(n_1_1_890), .A3(n_1_1_837), .A4(
      n_1_1_836), .ZN(n_1_1_835));
   AOI22_X1 i_1_1_850 (.A1(\mem[77] [13]), .A2(n_1_1_1133), .B1(n_1_1_1041), 
      .B2(\mem[7] [13]), .ZN(n_1_1_836));
   AOI22_X1 i_1_1_851 (.A1(\mem[0] [13]), .A2(n_1_1_1066), .B1(n_1_1_1049), 
      .B2(\mem[17] [13]), .ZN(n_1_1_837));
   NAND4_X1 i_1_1_852 (.A1(n_1_1_849), .A2(n_1_1_848), .A3(n_1_1_843), .A4(
      n_1_1_839), .ZN(n_1_1_838));
   AOI221_X1 i_1_1_853 (.A(n_1_1_840), .B1(n_1_1_1055), .B2(\mem[74] [13]), 
      .C1(\mem[76] [13]), .C2(n_1_1_1039), .ZN(n_1_1_839));
   NAND4_X1 i_1_1_854 (.A1(n_1_1_888), .A2(n_1_1_887), .A3(n_1_1_842), .A4(
      n_1_1_841), .ZN(n_1_1_840));
   AOI22_X1 i_1_1_855 (.A1(\mem[57] [13]), .A2(n_1_1_1108), .B1(n_1_1_1104), 
      .B2(\mem[48] [13]), .ZN(n_1_1_841));
   AOI22_X1 i_1_1_856 (.A1(\mem[79] [13]), .A2(n_1_1_1135), .B1(n_1_1_1073), 
      .B2(\mem[8] [13]), .ZN(n_1_1_842));
   AOI221_X1 i_1_1_857 (.A(n_1_1_844), .B1(n_1_1_1105), .B2(\mem[49] [13]), 
      .C1(\mem[51] [13]), .C2(n_1_1_1059), .ZN(n_1_1_843));
   NAND3_X1 i_1_1_858 (.A1(n_1_1_847), .A2(n_1_1_846), .A3(n_1_1_845), .ZN(
      n_1_1_844));
   AOI22_X1 i_1_1_859 (.A1(\mem[21] [13]), .A2(n_1_1_1081), .B1(n_1_1_1080), 
      .B2(\mem[19] [13]), .ZN(n_1_1_845));
   AOI22_X1 i_1_1_860 (.A1(\mem[54] [13]), .A2(n_1_1_1106), .B1(n_1_1_1030), 
      .B2(\mem[20] [13]), .ZN(n_1_1_846));
   AOI22_X1 i_1_1_861 (.A1(\mem[34] [13]), .A2(n_1_1_1093), .B1(n_1_1_1032), 
      .B2(\mem[44] [13]), .ZN(n_1_1_847));
   AOI22_X1 i_1_1_862 (.A1(\mem[59] [13]), .A2(n_1_1_1111), .B1(n_1_1_1025), 
      .B2(\mem[43] [13]), .ZN(n_1_1_848));
   AOI222_X1 i_1_1_863 (.A1(\mem[37] [13]), .A2(n_1_1_1096), .B1(n_1_1_1075), 
      .B2(\mem[13] [13]), .C1(n_1_1_1069), .C2(\mem[3] [13]), .ZN(n_1_1_849));
   NAND4_X1 i_1_1_864 (.A1(n_1_1_883), .A2(n_1_1_853), .A3(n_1_1_852), .A4(
      n_1_1_851), .ZN(n_1_1_850));
   AOI222_X1 i_1_1_865 (.A1(\mem[87] [13]), .A2(n_1_1_1144), .B1(n_1_1_1044), 
      .B2(\mem[26] [13]), .C1(n_1_1_1050), .C2(\mem[90] [13]), .ZN(n_1_1_851));
   AOI222_X1 i_1_1_866 (.A1(\mem[78] [13]), .A2(n_1_1_1134), .B1(n_1_1_1109), 
      .B2(\mem[58] [13]), .C1(n_1_1_1092), .C2(\mem[33] [13]), .ZN(n_1_1_852));
   AOI221_X1 i_1_1_867 (.A(n_1_1_854), .B1(n_1_1_1033), .B2(\mem[42] [13]), 
      .C1(\mem[65] [13]), .C2(n_1_1_1119), .ZN(n_1_1_853));
   NAND3_X1 i_1_1_868 (.A1(n_1_1_893), .A2(n_1_1_885), .A3(n_1_1_884), .ZN(
      n_1_1_854));
   AOI221_X1 i_1_1_869 (.A(n_1_1_856), .B1(n_1_1_1057), .B2(\mem[61] [13]), 
      .C1(\mem[94] [13]), .C2(n_1_1_1157), .ZN(n_1_1_855));
   NAND4_X1 i_1_1_870 (.A1(n_1_1_874), .A2(n_1_1_861), .A3(n_1_1_859), .A4(
      n_1_1_857), .ZN(n_1_1_856));
   AOI221_X1 i_1_1_871 (.A(n_1_1_858), .B1(n_1_1_1074), .B2(\mem[9] [13]), 
      .C1(\mem[31] [13]), .C2(n_1_1_1088), .ZN(n_1_1_857));
   NAND3_X1 i_1_1_872 (.A1(n_1_1_886), .A2(n_1_1_878), .A3(n_1_1_871), .ZN(
      n_1_1_858));
   AOI221_X1 i_1_1_873 (.A(n_1_1_860), .B1(n_1_1_1036), .B2(\mem[14] [13]), 
      .C1(\mem[68] [13]), .C2(n_1_1_1122), .ZN(n_1_1_859));
   NAND3_X1 i_1_1_874 (.A1(n_1_1_873), .A2(n_1_1_872), .A3(n_1_1_867), .ZN(
      n_1_1_860));
   NOR4_X1 i_1_1_875 (.A1(n_1_1_865), .A2(n_1_1_864), .A3(n_1_1_863), .A4(
      n_1_1_862), .ZN(n_1_1_861));
   NAND4_X1 i_1_1_876 (.A1(n_1_1_875), .A2(n_1_1_870), .A3(n_1_1_869), .A4(
      n_1_1_868), .ZN(n_1_1_862));
   NAND4_X1 i_1_1_877 (.A1(n_1_1_894), .A2(n_1_1_892), .A3(n_1_1_879), .A4(
      n_1_1_876), .ZN(n_1_1_863));
   NAND4_X1 i_1_1_878 (.A1(n_1_1_891), .A2(n_1_1_889), .A3(n_1_1_881), .A4(
      n_1_1_880), .ZN(n_1_1_864));
   NAND4_X1 i_1_1_879 (.A1(n_1_1_897), .A2(n_1_1_895), .A3(n_1_1_882), .A4(
      n_1_1_866), .ZN(n_1_1_865));
   AOI22_X1 i_1_1_880 (.A1(\mem[81] [13]), .A2(n_1_1_1139), .B1(n_1_1_1047), 
      .B2(\mem[83] [13]), .ZN(n_1_1_866));
   AOI22_X1 i_1_1_881 (.A1(\mem[41] [13]), .A2(n_1_1_1100), .B1(n_1_1_1048), 
      .B2(\mem[10] [13]), .ZN(n_1_1_867));
   AOI22_X1 i_1_1_882 (.A1(\mem[89] [13]), .A2(n_1_1_1148), .B1(n_1_1_1060), 
      .B2(\mem[28] [13]), .ZN(n_1_1_868));
   AOI22_X1 i_1_1_883 (.A1(\mem[84] [13]), .A2(n_1_1_1062), .B1(n_1_1_1056), 
      .B2(\mem[88] [13]), .ZN(n_1_1_869));
   AOI22_X1 i_1_1_884 (.A1(\mem[67] [13]), .A2(n_1_1_1121), .B1(n_1_1_1046), 
      .B2(\mem[60] [13]), .ZN(n_1_1_870));
   AOI22_X1 i_1_1_885 (.A1(\mem[70] [13]), .A2(n_1_1_1125), .B1(n_1_1_1068), 
      .B2(\mem[2] [13]), .ZN(n_1_1_871));
   AOI22_X1 i_1_1_886 (.A1(\mem[46] [13]), .A2(n_1_1_1101), .B1(n_1_1_1031), 
      .B2(\mem[39] [13]), .ZN(n_1_1_872));
   AOI22_X1 i_1_1_887 (.A1(\mem[40] [13]), .A2(n_1_1_1099), .B1(n_1_1_1070), 
      .B2(\mem[4] [13]), .ZN(n_1_1_873));
   AOI22_X1 i_1_1_888 (.A1(\mem[12] [13]), .A2(n_1_1_1042), .B1(n_1_1_1029), 
      .B2(\mem[62] [13]), .ZN(n_1_1_874));
   AOI22_X1 i_1_1_889 (.A1(\mem[93] [13]), .A2(n_1_1_1155), .B1(n_1_1_1028), 
      .B2(\mem[82] [13]), .ZN(n_1_1_875));
   AOI22_X1 i_1_1_890 (.A1(\mem[71] [13]), .A2(n_1_1_1126), .B1(n_1_1_1083), 
      .B2(\mem[24] [13]), .ZN(n_1_1_876));
   AOI22_X1 i_1_1_891 (.A1(\mem[32] [13]), .A2(n_1_1_1091), .B1(n_1_1_1052), 
      .B2(\mem[23] [13]), .ZN(n_1_1_877));
   AOI22_X1 i_1_1_892 (.A1(\mem[73] [13]), .A2(n_1_1_1129), .B1(n_1_1_1118), 
      .B2(\mem[64] [13]), .ZN(n_1_1_878));
   AOI22_X1 i_1_1_893 (.A1(\mem[80] [13]), .A2(n_1_1_1138), .B1(n_1_1_1095), 
      .B2(\mem[36] [13]), .ZN(n_1_1_879));
   AOI22_X1 i_1_1_894 (.A1(\mem[75] [13]), .A2(n_1_1_1061), .B1(n_1_1_1035), 
      .B2(\mem[50] [13]), .ZN(n_1_1_880));
   AOI22_X1 i_1_1_895 (.A1(\mem[96] [13]), .A2(n_1_1_1163), .B1(n_1_1_1051), 
      .B2(\mem[29] [13]), .ZN(n_1_1_881));
   AOI22_X1 i_1_1_896 (.A1(\mem[5] [13]), .A2(n_1_1_1071), .B1(n_1_1_1063), 
      .B2(\mem[11] [13]), .ZN(n_1_1_882));
   AOI22_X1 i_1_1_897 (.A1(\mem[30] [13]), .A2(n_1_1_1087), .B1(n_1_1_1037), 
      .B2(\mem[91] [13]), .ZN(n_1_1_883));
   AOI22_X1 i_1_1_898 (.A1(\mem[45] [13]), .A2(n_1_1_1045), .B1(n_1_1_1040), 
      .B2(\mem[52] [13]), .ZN(n_1_1_884));
   AOI22_X1 i_1_1_899 (.A1(\mem[86] [13]), .A2(n_1_1_1142), .B1(n_1_1_1038), 
      .B2(\mem[15] [13]), .ZN(n_1_1_885));
   AOI22_X1 i_1_1_900 (.A1(\mem[66] [13]), .A2(n_1_1_1120), .B1(n_1_1_1064), 
      .B2(\mem[18] [13]), .ZN(n_1_1_886));
   AOI22_X1 i_1_1_901 (.A1(\mem[98] [13]), .A2(n_1_1_1168), .B1(n_1_1_1107), 
      .B2(\mem[55] [13]), .ZN(n_1_1_887));
   AOI22_X1 i_1_1_902 (.A1(\mem[92] [13]), .A2(n_1_1_1153), .B1(n_1_1_1054), 
      .B2(\mem[22] [13]), .ZN(n_1_1_888));
   AOI22_X1 i_1_1_903 (.A1(\mem[47] [13]), .A2(n_1_1_1102), .B1(n_1_1_1053), 
      .B2(\mem[95] [13]), .ZN(n_1_1_889));
   AOI22_X1 i_1_1_904 (.A1(\mem[6] [13]), .A2(n_1_1_1072), .B1(n_1_1_1027), 
      .B2(\mem[27] [13]), .ZN(n_1_1_890));
   AOI22_X1 i_1_1_905 (.A1(\mem[97] [13]), .A2(n_1_1_1165), .B1(n_1_1_1116), 
      .B2(\mem[63] [13]), .ZN(n_1_1_891));
   AOI22_X1 i_1_1_906 (.A1(\mem[35] [13]), .A2(n_1_1_1094), .B1(n_1_1_1026), 
      .B2(\mem[56] [13]), .ZN(n_1_1_892));
   AOI22_X1 i_1_1_907 (.A1(\mem[25] [13]), .A2(n_1_1_1084), .B1(n_1_1_1078), 
      .B2(\mem[16] [13]), .ZN(n_1_1_893));
   AOI22_X1 i_1_1_908 (.A1(\mem[69] [13]), .A2(n_1_1_1123), .B1(n_1_1_1043), 
      .B2(\mem[53] [13]), .ZN(n_1_1_894));
   AOI22_X1 i_1_1_909 (.A1(\mem[100] [13]), .A2(n_1_1_1174), .B1(n_1_1_1067), 
      .B2(\mem[1] [13]), .ZN(n_1_1_895));
   AOI22_X1 i_1_1_910 (.A1(\mem[99] [13]), .A2(n_1_1_1171), .B1(n_1_1_1127), 
      .B2(\mem[72] [13]), .ZN(n_1_1_896));
   AOI22_X1 i_1_1_911 (.A1(\mem[38] [13]), .A2(n_1_1_1097), .B1(n_1_1_1058), 
      .B2(\mem[85] [13]), .ZN(n_1_1_897));
   AOI21_X1 i_1_1_912 (.A(n_1_1_963), .B1(n_1_1_898), .B2(read_signal), .ZN(
      n_1_14));
   NOR3_X1 i_1_1_913 (.A1(n_1_1_920), .A2(n_1_1_914), .A3(n_1_1_899), .ZN(
      n_1_1_898));
   NAND4_X1 i_1_1_914 (.A1(n_1_1_954), .A2(n_1_1_904), .A3(n_1_1_903), .A4(
      n_1_1_900), .ZN(n_1_1_899));
   AOI221_X1 i_1_1_915 (.A(n_1_1_901), .B1(n_1_1_1052), .B2(\mem[23] [14]), 
      .C1(\mem[94] [14]), .C2(n_1_1_1157), .ZN(n_1_1_900));
   NAND4_X1 i_1_1_916 (.A1(n_1_1_955), .A2(n_1_1_953), .A3(n_1_1_952), .A4(
      n_1_1_902), .ZN(n_1_1_901));
   AOI22_X1 i_1_1_917 (.A1(\mem[32] [14]), .A2(n_1_1_1091), .B1(n_1_1_1045), 
      .B2(\mem[45] [14]), .ZN(n_1_1_902));
   AOI22_X1 i_1_1_918 (.A1(\mem[79] [14]), .A2(n_1_1_1135), .B1(n_1_1_1078), 
      .B2(\mem[16] [14]), .ZN(n_1_1_903));
   NOR4_X1 i_1_1_919 (.A1(n_1_1_911), .A2(n_1_1_909), .A3(n_1_1_907), .A4(
      n_1_1_905), .ZN(n_1_1_904));
   NAND4_X1 i_1_1_920 (.A1(n_1_1_956), .A2(n_1_1_944), .A3(n_1_1_943), .A4(
      n_1_1_906), .ZN(n_1_1_905));
   AOI22_X1 i_1_1_921 (.A1(\mem[87] [14]), .A2(n_1_1_1144), .B1(n_1_1_1044), 
      .B2(\mem[26] [14]), .ZN(n_1_1_906));
   NAND4_X1 i_1_1_922 (.A1(n_1_1_961), .A2(n_1_1_950), .A3(n_1_1_949), .A4(
      n_1_1_908), .ZN(n_1_1_907));
   AOI22_X1 i_1_1_923 (.A1(\mem[5] [14]), .A2(n_1_1_1071), .B1(n_1_1_1029), 
      .B2(\mem[62] [14]), .ZN(n_1_1_908));
   NAND4_X1 i_1_1_924 (.A1(n_1_1_948), .A2(n_1_1_942), .A3(n_1_1_941), .A4(
      n_1_1_910), .ZN(n_1_1_909));
   AOI22_X1 i_1_1_925 (.A1(\mem[46] [14]), .A2(n_1_1_1101), .B1(n_1_1_1036), 
      .B2(\mem[14] [14]), .ZN(n_1_1_910));
   NAND4_X1 i_1_1_926 (.A1(n_1_1_958), .A2(n_1_1_951), .A3(n_1_1_913), .A4(
      n_1_1_912), .ZN(n_1_1_911));
   AOI22_X1 i_1_1_927 (.A1(\mem[4] [14]), .A2(n_1_1_1070), .B1(n_1_1_1062), 
      .B2(\mem[84] [14]), .ZN(n_1_1_912));
   AOI22_X1 i_1_1_928 (.A1(\mem[98] [14]), .A2(n_1_1_1168), .B1(n_1_1_1054), 
      .B2(\mem[22] [14]), .ZN(n_1_1_913));
   NAND4_X1 i_1_1_929 (.A1(n_1_1_919), .A2(n_1_1_918), .A3(n_1_1_917), .A4(
      n_1_1_915), .ZN(n_1_1_914));
   AOI221_X1 i_1_1_930 (.A(n_1_1_916), .B1(n_1_1_1099), .B2(\mem[40] [14]), 
      .C1(\mem[99] [14]), .C2(n_1_1_1171), .ZN(n_1_1_915));
   NAND3_X1 i_1_1_931 (.A1(n_1_1_959), .A2(n_1_1_939), .A3(n_1_1_938), .ZN(
      n_1_1_916));
   AOI222_X1 i_1_1_932 (.A1(\mem[95] [14]), .A2(n_1_1_1053), .B1(n_1_1_1046), 
      .B2(\mem[60] [14]), .C1(n_1_1_1038), .C2(\mem[15] [14]), .ZN(n_1_1_917));
   AOI22_X1 i_1_1_933 (.A1(\mem[96] [14]), .A2(n_1_1_1163), .B1(n_1_1_1094), 
      .B2(\mem[35] [14]), .ZN(n_1_1_918));
   AOI22_X1 i_1_1_934 (.A1(\mem[66] [14]), .A2(n_1_1_1120), .B1(n_1_1_1109), 
      .B2(\mem[58] [14]), .ZN(n_1_1_919));
   NAND4_X1 i_1_1_935 (.A1(n_1_1_940), .A2(n_1_1_937), .A3(n_1_1_936), .A4(
      n_1_1_921), .ZN(n_1_1_920));
   AOI211_X1 i_1_1_936 (.A(n_1_1_932), .B(n_1_1_922), .C1(\mem[17] [14]), 
      .C2(n_1_1_1049), .ZN(n_1_1_921));
   NAND3_X1 i_1_1_937 (.A1(n_1_1_929), .A2(n_1_1_927), .A3(n_1_1_923), .ZN(
      n_1_1_922));
   AOI221_X1 i_1_1_938 (.A(n_1_1_924), .B1(n_1_1_1063), .B2(\mem[11] [14]), 
      .C1(\mem[25] [14]), .C2(n_1_1_1084), .ZN(n_1_1_923));
   NAND3_X1 i_1_1_939 (.A1(n_1_1_945), .A2(n_1_1_926), .A3(n_1_1_925), .ZN(
      n_1_1_924));
   AOI22_X1 i_1_1_940 (.A1(\mem[51] [14]), .A2(n_1_1_1059), .B1(n_1_1_1050), 
      .B2(\mem[90] [14]), .ZN(n_1_1_925));
   AOI22_X1 i_1_1_941 (.A1(\mem[38] [14]), .A2(n_1_1_1097), .B1(n_1_1_1066), 
      .B2(\mem[0] [14]), .ZN(n_1_1_926));
   AOI221_X1 i_1_1_942 (.A(n_1_1_928), .B1(n_1_1_1068), .B2(\mem[2] [14]), 
      .C1(\mem[61] [14]), .C2(n_1_1_1057), .ZN(n_1_1_927));
   NAND3_X1 i_1_1_943 (.A1(n_1_1_960), .A2(n_1_1_947), .A3(n_1_1_946), .ZN(
      n_1_1_928));
   AOI221_X1 i_1_1_944 (.A(n_1_1_930), .B1(n_1_1_1055), .B2(\mem[74] [14]), 
      .C1(\mem[86] [14]), .C2(n_1_1_1142), .ZN(n_1_1_929));
   NAND3_X1 i_1_1_945 (.A1(n_1_1_962), .A2(n_1_1_957), .A3(n_1_1_931), .ZN(
      n_1_1_930));
   AOI22_X1 i_1_1_946 (.A1(\mem[55] [14]), .A2(n_1_1_1107), .B1(n_1_1_1048), 
      .B2(\mem[10] [14]), .ZN(n_1_1_931));
   NAND3_X1 i_1_1_947 (.A1(n_1_1_935), .A2(n_1_1_934), .A3(n_1_1_933), .ZN(
      n_1_1_932));
   AOI222_X1 i_1_1_948 (.A1(\mem[57] [14]), .A2(n_1_1_1108), .B1(n_1_1_1083), 
      .B2(\mem[24] [14]), .C1(n_1_1_1039), .C2(\mem[76] [14]), .ZN(n_1_1_933));
   AOI22_X1 i_1_1_949 (.A1(\mem[67] [14]), .A2(n_1_1_1121), .B1(n_1_1_1058), 
      .B2(\mem[85] [14]), .ZN(n_1_1_934));
   AOI22_X1 i_1_1_950 (.A1(\mem[92] [14]), .A2(n_1_1_1153), .B1(n_1_1_1067), 
      .B2(\mem[1] [14]), .ZN(n_1_1_935));
   AOI22_X1 i_1_1_951 (.A1(\mem[44] [14]), .A2(n_1_1_1032), .B1(n_1_1_1030), 
      .B2(\mem[20] [14]), .ZN(n_1_1_936));
   AOI222_X1 i_1_1_952 (.A1(\mem[37] [14]), .A2(n_1_1_1096), .B1(n_1_1_1088), 
      .B2(\mem[31] [14]), .C1(n_1_1_1060), .C2(\mem[28] [14]), .ZN(n_1_1_937));
   AOI22_X1 i_1_1_953 (.A1(\mem[49] [14]), .A2(n_1_1_1105), .B1(n_1_1_1061), 
      .B2(\mem[75] [14]), .ZN(n_1_1_938));
   AOI22_X1 i_1_1_954 (.A1(\mem[93] [14]), .A2(n_1_1_1155), .B1(n_1_1_1028), 
      .B2(\mem[82] [14]), .ZN(n_1_1_939));
   AOI222_X1 i_1_1_955 (.A1(\mem[97] [14]), .A2(n_1_1_1165), .B1(n_1_1_1138), 
      .B2(\mem[80] [14]), .C1(n_1_1_1126), .C2(\mem[71] [14]), .ZN(n_1_1_940));
   AOI22_X1 i_1_1_956 (.A1(\mem[63] [14]), .A2(n_1_1_1116), .B1(n_1_1_1026), 
      .B2(\mem[56] [14]), .ZN(n_1_1_941));
   AOI22_X1 i_1_1_957 (.A1(\mem[65] [14]), .A2(n_1_1_1119), .B1(n_1_1_1043), 
      .B2(\mem[53] [14]), .ZN(n_1_1_942));
   AOI22_X1 i_1_1_958 (.A1(\mem[100] [14]), .A2(n_1_1_1174), .B1(n_1_1_1042), 
      .B2(\mem[12] [14]), .ZN(n_1_1_943));
   AOI22_X1 i_1_1_959 (.A1(\mem[30] [14]), .A2(n_1_1_1087), .B1(n_1_1_1047), 
      .B2(\mem[83] [14]), .ZN(n_1_1_944));
   AOI22_X1 i_1_1_960 (.A1(\mem[68] [14]), .A2(n_1_1_1122), .B1(n_1_1_1075), 
      .B2(\mem[13] [14]), .ZN(n_1_1_945));
   AOI22_X1 i_1_1_961 (.A1(\mem[72] [14]), .A2(n_1_1_1127), .B1(n_1_1_1073), 
      .B2(\mem[8] [14]), .ZN(n_1_1_946));
   AOI22_X1 i_1_1_962 (.A1(\mem[47] [14]), .A2(n_1_1_1102), .B1(n_1_1_1041), 
      .B2(\mem[7] [14]), .ZN(n_1_1_947));
   AOI22_X1 i_1_1_963 (.A1(\mem[21] [14]), .A2(n_1_1_1081), .B1(n_1_1_1031), 
      .B2(\mem[39] [14]), .ZN(n_1_1_948));
   AOI22_X1 i_1_1_964 (.A1(\mem[64] [14]), .A2(n_1_1_1118), .B1(n_1_1_1064), 
      .B2(\mem[18] [14]), .ZN(n_1_1_949));
   AOI22_X1 i_1_1_965 (.A1(\mem[54] [14]), .A2(n_1_1_1106), .B1(n_1_1_1025), 
      .B2(\mem[43] [14]), .ZN(n_1_1_950));
   AOI22_X1 i_1_1_966 (.A1(\mem[89] [14]), .A2(n_1_1_1148), .B1(n_1_1_1072), 
      .B2(\mem[6] [14]), .ZN(n_1_1_951));
   AOI22_X1 i_1_1_967 (.A1(\mem[3] [14]), .A2(n_1_1_1069), .B1(n_1_1_1040), 
      .B2(\mem[52] [14]), .ZN(n_1_1_952));
   AOI22_X1 i_1_1_968 (.A1(\mem[41] [14]), .A2(n_1_1_1100), .B1(n_1_1_1051), 
      .B2(\mem[29] [14]), .ZN(n_1_1_953));
   AOI22_X1 i_1_1_969 (.A1(\mem[78] [14]), .A2(n_1_1_1134), .B1(n_1_1_1033), 
      .B2(\mem[42] [14]), .ZN(n_1_1_954));
   AOI22_X1 i_1_1_970 (.A1(\mem[48] [14]), .A2(n_1_1_1104), .B1(n_1_1_1035), 
      .B2(\mem[50] [14]), .ZN(n_1_1_955));
   AOI22_X1 i_1_1_971 (.A1(\mem[73] [14]), .A2(n_1_1_1129), .B1(n_1_1_1080), 
      .B2(\mem[19] [14]), .ZN(n_1_1_956));
   AOI22_X1 i_1_1_972 (.A1(\mem[70] [14]), .A2(n_1_1_1125), .B1(n_1_1_1092), 
      .B2(\mem[33] [14]), .ZN(n_1_1_957));
   AOI22_X1 i_1_1_973 (.A1(\mem[81] [14]), .A2(n_1_1_1139), .B1(n_1_1_1056), 
      .B2(\mem[88] [14]), .ZN(n_1_1_958));
   AOI22_X1 i_1_1_974 (.A1(\mem[77] [14]), .A2(n_1_1_1133), .B1(n_1_1_1123), 
      .B2(\mem[69] [14]), .ZN(n_1_1_959));
   AOI22_X1 i_1_1_975 (.A1(\mem[59] [14]), .A2(n_1_1_1111), .B1(n_1_1_1027), 
      .B2(\mem[27] [14]), .ZN(n_1_1_960));
   AOI22_X1 i_1_1_976 (.A1(\mem[34] [14]), .A2(n_1_1_1093), .B1(n_1_1_1074), 
      .B2(\mem[9] [14]), .ZN(n_1_1_961));
   AOI22_X1 i_1_1_977 (.A1(\mem[36] [14]), .A2(n_1_1_1095), .B1(n_1_1_1037), 
      .B2(\mem[91] [14]), .ZN(n_1_1_962));
   NOR2_X1 i_1_1_978 (.A1(read_signal), .A2(dataout[14]), .ZN(n_1_1_963));
   MUX2_X1 i_1_1_979 (.A(dataout[15]), .B(n_1_1_964), .S(read_signal), .Z(n_1_15));
   NAND4_X1 i_1_1_980 (.A1(n_1_1_1017), .A2(n_1_1_1011), .A3(n_1_1_1005), 
      .A4(n_1_1_965), .ZN(n_1_1_964));
   AOI221_X1 i_1_1_981 (.A(n_1_1_966), .B1(n_1_1_1100), .B2(\mem[41] [15]), 
      .C1(\mem[42] [15]), .C2(n_1_1_1033), .ZN(n_1_1_965));
   NAND4_X1 i_1_1_982 (.A1(n_1_1_997), .A2(n_1_1_991), .A3(n_1_1_972), .A4(
      n_1_1_967), .ZN(n_1_1_966));
   AOI221_X1 i_1_1_983 (.A(n_1_1_968), .B1(n_1_1_1031), .B2(\mem[39] [15]), 
      .C1(\mem[62] [15]), .C2(n_1_1_1029), .ZN(n_1_1_967));
   NAND3_X1 i_1_1_984 (.A1(n_1_1_971), .A2(n_1_1_970), .A3(n_1_1_969), .ZN(
      n_1_1_968));
   AOI22_X1 i_1_1_985 (.A1(\mem[21] [15]), .A2(n_1_1_1081), .B1(n_1_1_1060), 
      .B2(\mem[28] [15]), .ZN(n_1_1_969));
   AOI22_X1 i_1_1_986 (.A1(\mem[57] [15]), .A2(n_1_1_1108), .B1(n_1_1_1080), 
      .B2(\mem[19] [15]), .ZN(n_1_1_970));
   AOI22_X1 i_1_1_987 (.A1(\mem[75] [15]), .A2(n_1_1_1061), .B1(n_1_1_1042), 
      .B2(\mem[12] [15]), .ZN(n_1_1_971));
   NOR4_X1 i_1_1_988 (.A1(n_1_1_987), .A2(n_1_1_982), .A3(n_1_1_978), .A4(
      n_1_1_973), .ZN(n_1_1_972));
   NAND4_X1 i_1_1_989 (.A1(n_1_1_977), .A2(n_1_1_976), .A3(n_1_1_975), .A4(
      n_1_1_974), .ZN(n_1_1_973));
   AOI22_X1 i_1_1_990 (.A1(\mem[96] [15]), .A2(n_1_1_1163), .B1(n_1_1_1101), 
      .B2(\mem[46] [15]), .ZN(n_1_1_974));
   AOI22_X1 i_1_1_991 (.A1(\mem[69] [15]), .A2(n_1_1_1123), .B1(n_1_1_1096), 
      .B2(\mem[37] [15]), .ZN(n_1_1_975));
   AOI22_X1 i_1_1_992 (.A1(\mem[52] [15]), .A2(n_1_1_1040), .B1(n_1_1_1030), 
      .B2(\mem[20] [15]), .ZN(n_1_1_976));
   AOI22_X1 i_1_1_993 (.A1(\mem[66] [15]), .A2(n_1_1_1120), .B1(n_1_1_1105), 
      .B2(\mem[49] [15]), .ZN(n_1_1_977));
   NAND4_X1 i_1_1_994 (.A1(n_1_1_1024), .A2(n_1_1_981), .A3(n_1_1_980), .A4(
      n_1_1_979), .ZN(n_1_1_978));
   AOI22_X1 i_1_1_995 (.A1(\mem[92] [15]), .A2(n_1_1_1153), .B1(n_1_1_1072), 
      .B2(\mem[6] [15]), .ZN(n_1_1_979));
   AOI22_X1 i_1_1_996 (.A1(\mem[87] [15]), .A2(n_1_1_1144), .B1(n_1_1_1083), 
      .B2(\mem[24] [15]), .ZN(n_1_1_980));
   AOI22_X1 i_1_1_997 (.A1(\mem[98] [15]), .A2(n_1_1_1168), .B1(n_1_1_1056), 
      .B2(\mem[88] [15]), .ZN(n_1_1_981));
   NAND4_X1 i_1_1_998 (.A1(n_1_1_986), .A2(n_1_1_985), .A3(n_1_1_984), .A4(
      n_1_1_983), .ZN(n_1_1_982));
   AOI22_X1 i_1_1_999 (.A1(\mem[99] [15]), .A2(n_1_1_1171), .B1(n_1_1_1078), 
      .B2(\mem[16] [15]), .ZN(n_1_1_983));
   AOI22_X1 i_1_1_1000 (.A1(\mem[72] [15]), .A2(n_1_1_1127), .B1(n_1_1_1043), 
      .B2(\mem[53] [15]), .ZN(n_1_1_984));
   AOI22_X1 i_1_1_1001 (.A1(\mem[44] [15]), .A2(n_1_1_1032), .B1(n_1_1_1025), 
      .B2(\mem[43] [15]), .ZN(n_1_1_985));
   AOI22_X1 i_1_1_1002 (.A1(\mem[100] [15]), .A2(n_1_1_1174), .B1(n_1_1_1058), 
      .B2(\mem[85] [15]), .ZN(n_1_1_986));
   NAND3_X1 i_1_1_1003 (.A1(n_1_1_990), .A2(n_1_1_989), .A3(n_1_1_988), .ZN(
      n_1_1_987));
   AOI22_X1 i_1_1_1004 (.A1(\mem[25] [15]), .A2(n_1_1_1084), .B1(n_1_1_1044), 
      .B2(\mem[26] [15]), .ZN(n_1_1_988));
   AOI222_X1 i_1_1_1005 (.A1(\mem[73] [15]), .A2(n_1_1_1129), .B1(n_1_1_1057), 
      .B2(\mem[61] [15]), .C1(n_1_1_1050), .C2(\mem[90] [15]), .ZN(n_1_1_989));
   AOI222_X1 i_1_1_1006 (.A1(\mem[81] [15]), .A2(n_1_1_1139), .B1(n_1_1_1055), 
      .B2(\mem[74] [15]), .C1(n_1_1_1054), .C2(\mem[22] [15]), .ZN(n_1_1_990));
   AOI221_X1 i_1_1_1007 (.A(n_1_1_992), .B1(n_1_1_1027), .B2(\mem[27] [15]), 
      .C1(\mem[82] [15]), .C2(n_1_1_1028), .ZN(n_1_1_991));
   NAND4_X1 i_1_1_1008 (.A1(n_1_1_996), .A2(n_1_1_995), .A3(n_1_1_994), .A4(
      n_1_1_993), .ZN(n_1_1_992));
   AOI22_X1 i_1_1_1009 (.A1(\mem[51] [15]), .A2(n_1_1_1059), .B1(n_1_1_1045), 
      .B2(\mem[45] [15]), .ZN(n_1_1_993));
   AOI22_X1 i_1_1_1010 (.A1(\mem[67] [15]), .A2(n_1_1_1121), .B1(n_1_1_1046), 
      .B2(\mem[60] [15]), .ZN(n_1_1_994));
   AOI22_X1 i_1_1_1011 (.A1(\mem[54] [15]), .A2(n_1_1_1106), .B1(n_1_1_1039), 
      .B2(\mem[76] [15]), .ZN(n_1_1_995));
   AOI22_X1 i_1_1_1012 (.A1(\mem[79] [15]), .A2(n_1_1_1135), .B1(n_1_1_1053), 
      .B2(\mem[95] [15]), .ZN(n_1_1_996));
   AOI221_X1 i_1_1_1013 (.A(n_1_1_998), .B1(n_1_1_1049), .B2(\mem[17] [15]), 
      .C1(\mem[30] [15]), .C2(n_1_1_1087), .ZN(n_1_1_997));
   NAND3_X1 i_1_1_1014 (.A1(n_1_1_1001), .A2(n_1_1_1000), .A3(n_1_1_999), 
      .ZN(n_1_1_998));
   AOI222_X1 i_1_1_1015 (.A1(\mem[68] [15]), .A2(n_1_1_1122), .B1(n_1_1_1075), 
      .B2(\mem[13] [15]), .C1(n_1_1_1064), .C2(\mem[18] [15]), .ZN(n_1_1_999));
   AOI222_X1 i_1_1_1016 (.A1(\mem[89] [15]), .A2(n_1_1_1148), .B1(n_1_1_1097), 
      .B2(\mem[38] [15]), .C1(n_1_1_1066), .C2(\mem[0] [15]), .ZN(n_1_1_1000));
   AOI221_X1 i_1_1_1017 (.A(n_1_1_1002), .B1(n_1_1_1036), .B2(\mem[14] [15]), 
      .C1(\mem[55] [15]), .C2(n_1_1_1107), .ZN(n_1_1_1001));
   NAND3_X1 i_1_1_1018 (.A1(n_1_1_1065), .A2(n_1_1_1004), .A3(n_1_1_1003), 
      .ZN(n_1_1_1002));
   AOI22_X1 i_1_1_1019 (.A1(\mem[47] [15]), .A2(n_1_1_1102), .B1(n_1_1_1052), 
      .B2(\mem[23] [15]), .ZN(n_1_1_1003));
   AOI22_X1 i_1_1_1020 (.A1(\mem[4] [15]), .A2(n_1_1_1070), .B1(n_1_1_1048), 
      .B2(\mem[10] [15]), .ZN(n_1_1_1004));
   AOI221_X1 i_1_1_1021 (.A(n_1_1_1006), .B1(n_1_1_1041), .B2(\mem[7] [15]), 
      .C1(\mem[97] [15]), .C2(n_1_1_1165), .ZN(n_1_1_1005));
   NAND4_X1 i_1_1_1022 (.A1(n_1_1_1010), .A2(n_1_1_1009), .A3(n_1_1_1008), 
      .A4(n_1_1_1007), .ZN(n_1_1_1006));
   AOI22_X1 i_1_1_1023 (.A1(\mem[64] [15]), .A2(n_1_1_1118), .B1(n_1_1_1067), 
      .B2(\mem[1] [15]), .ZN(n_1_1_1007));
   AOI22_X1 i_1_1_1024 (.A1(\mem[78] [15]), .A2(n_1_1_1134), .B1(n_1_1_1069), 
      .B2(\mem[3] [15]), .ZN(n_1_1_1008));
   AOI22_X1 i_1_1_1025 (.A1(\mem[93] [15]), .A2(n_1_1_1155), .B1(n_1_1_1109), 
      .B2(\mem[58] [15]), .ZN(n_1_1_1009));
   AOI22_X1 i_1_1_1026 (.A1(\mem[34] [15]), .A2(n_1_1_1093), .B1(n_1_1_1047), 
      .B2(\mem[83] [15]), .ZN(n_1_1_1010));
   AOI221_X1 i_1_1_1027 (.A(n_1_1_1012), .B1(n_1_1_1038), .B2(\mem[15] [15]), 
      .C1(\mem[91] [15]), .C2(n_1_1_1037), .ZN(n_1_1_1011));
   NAND3_X1 i_1_1_1028 (.A1(n_1_1_1015), .A2(n_1_1_1014), .A3(n_1_1_1013), 
      .ZN(n_1_1_1012));
   AOI22_X1 i_1_1_1029 (.A1(\mem[70] [15]), .A2(n_1_1_1125), .B1(n_1_1_1111), 
      .B2(\mem[59] [15]), .ZN(n_1_1_1013));
   AOI222_X1 i_1_1_1030 (.A1(\mem[80] [15]), .A2(n_1_1_1138), .B1(n_1_1_1104), 
      .B2(\mem[48] [15]), .C1(n_1_1_1094), .C2(\mem[35] [15]), .ZN(n_1_1_1014));
   AOI221_X1 i_1_1_1031 (.A(n_1_1_1016), .B1(n_1_1_1071), .B2(\mem[5] [15]), 
      .C1(\mem[8] [15]), .C2(n_1_1_1073), .ZN(n_1_1_1015));
   NAND3_X1 i_1_1_1032 (.A1(n_1_1_1020), .A2(n_1_1_1019), .A3(n_1_1_1018), 
      .ZN(n_1_1_1016));
   AOI221_X1 i_1_1_1033 (.A(n_1_1_1021), .B1(n_1_1_1051), .B2(\mem[29] [15]), 
      .C1(\mem[71] [15]), .C2(n_1_1_1126), .ZN(n_1_1_1017));
   AOI22_X1 i_1_1_1034 (.A1(\mem[94] [15]), .A2(n_1_1_1157), .B1(n_1_1_1133), 
      .B2(\mem[77] [15]), .ZN(n_1_1_1018));
   AOI22_X1 i_1_1_1035 (.A1(\mem[65] [15]), .A2(n_1_1_1119), .B1(n_1_1_1068), 
      .B2(\mem[2] [15]), .ZN(n_1_1_1019));
   AOI22_X1 i_1_1_1036 (.A1(\mem[86] [15]), .A2(n_1_1_1142), .B1(n_1_1_1088), 
      .B2(\mem[31] [15]), .ZN(n_1_1_1020));
   NAND3_X1 i_1_1_1037 (.A1(n_1_1_1034), .A2(n_1_1_1023), .A3(n_1_1_1022), 
      .ZN(n_1_1_1021));
   AOI22_X1 i_1_1_1038 (.A1(\mem[11] [15]), .A2(n_1_1_1063), .B1(n_1_1_1026), 
      .B2(\mem[56] [15]), .ZN(n_1_1_1022));
   AOI22_X1 i_1_1_1039 (.A1(\mem[32] [15]), .A2(n_1_1_1091), .B1(n_1_1_1062), 
      .B2(\mem[84] [15]), .ZN(n_1_1_1023));
   AOI22_X1 i_1_1_1040 (.A1(\mem[40] [15]), .A2(n_1_1_1099), .B1(n_1_1_1092), 
      .B2(\mem[33] [15]), .ZN(n_1_1_1024));
   NOR2_X1 i_1_1_1041 (.A1(n_1_1_1112), .A2(n_1_1_1103), .ZN(n_1_1_1025));
   NOR2_X1 i_1_1_1042 (.A1(n_1_1_1128), .A2(n_1_1_1117), .ZN(n_1_1_1026));
   NOR2_X1 i_1_1_1043 (.A1(n_1_1_1112), .A2(n_1_1_1089), .ZN(n_1_1_1027));
   NOR2_X1 i_1_1_1044 (.A1(n_1_1_1169), .A2(n_1_1_1159), .ZN(n_1_1_1028));
   NOR2_X1 i_1_1_1045 (.A1(n_1_1_1158), .A2(n_1_1_1117), .ZN(n_1_1_1029));
   NOR2_X1 i_1_1_1046 (.A1(n_1_1_1176), .A2(n_1_1_1089), .ZN(n_1_1_1030));
   NOR2_X1 i_1_1_1047 (.A1(n_1_1_1145), .A2(n_1_1_1103), .ZN(n_1_1_1031));
   NOR2_X1 i_1_1_1048 (.A1(n_1_1_1154), .A2(n_1_1_1103), .ZN(n_1_1_1032));
   NOR2_X1 i_1_1_1049 (.A1(n_1_1_1110), .A2(n_1_1_1103), .ZN(n_1_1_1033));
   AOI22_X1 i_1_1_1050 (.A1(\mem[36] [15]), .A2(n_1_1_1095), .B1(n_1_1_1035), 
      .B2(\mem[50] [15]), .ZN(n_1_1_1034));
   NOR2_X1 i_1_1_1051 (.A1(n_1_1_1169), .A2(n_1_1_1117), .ZN(n_1_1_1035));
   NOR2_X1 i_1_1_1052 (.A1(n_1_1_1158), .A2(n_1_1_1076), .ZN(n_1_1_1036));
   NOR2_X1 i_1_1_1053 (.A1(n_1_1_1159), .A2(n_1_1_1112), .ZN(n_1_1_1037));
   NOR2_X1 i_1_1_1054 (.A1(n_1_1_1137), .A2(n_1_1_1076), .ZN(n_1_1_1038));
   NOR2_X1 i_1_1_1055 (.A1(n_1_1_1154), .A2(n_1_1_1136), .ZN(n_1_1_1039));
   NOR2_X1 i_1_1_1056 (.A1(n_1_1_1176), .A2(n_1_1_1117), .ZN(n_1_1_1040));
   NOR2_X1 i_1_1_1057 (.A1(n_1_1_1145), .A2(n_1_1_1076), .ZN(n_1_1_1041));
   NOR2_X1 i_1_1_1058 (.A1(n_1_1_1154), .A2(n_1_1_1076), .ZN(n_1_1_1042));
   NOR2_X1 i_1_1_1059 (.A1(n_1_1_1124), .A2(n_1_1_1117), .ZN(n_1_1_1043));
   NOR2_X1 i_1_1_1060 (.A1(n_1_1_1110), .A2(n_1_1_1089), .ZN(n_1_1_1044));
   NOR2_X1 i_1_1_1061 (.A1(n_1_1_1156), .A2(n_1_1_1103), .ZN(n_1_1_1045));
   NOR2_X1 i_1_1_1062 (.A1(n_1_1_1154), .A2(n_1_1_1117), .ZN(n_1_1_1046));
   NOR2_X1 i_1_1_1063 (.A1(n_1_1_1172), .A2(n_1_1_1159), .ZN(n_1_1_1047));
   NOR2_X1 i_1_1_1064 (.A1(n_1_1_1110), .A2(n_1_1_1076), .ZN(n_1_1_1048));
   NOR2_X1 i_1_1_1065 (.A1(n_1_1_1166), .A2(n_1_1_1089), .ZN(n_1_1_1049));
   NOR2_X1 i_1_1_1066 (.A1(n_1_1_1159), .A2(n_1_1_1110), .ZN(n_1_1_1050));
   NOR2_X1 i_1_1_1067 (.A1(n_1_1_1156), .A2(n_1_1_1089), .ZN(n_1_1_1051));
   NOR2_X1 i_1_1_1068 (.A1(n_1_1_1145), .A2(n_1_1_1089), .ZN(n_1_1_1052));
   NOR2_X1 i_1_1_1069 (.A1(n_1_1_1159), .A2(n_1_1_1137), .ZN(n_1_1_1053));
   NOR2_X1 i_1_1_1070 (.A1(n_1_1_1143), .A2(n_1_1_1089), .ZN(n_1_1_1054));
   NOR2_X1 i_1_1_1071 (.A1(n_1_1_1136), .A2(n_1_1_1110), .ZN(n_1_1_1055));
   NOR2_X1 i_1_1_1072 (.A1(n_1_1_1159), .A2(n_1_1_1128), .ZN(n_1_1_1056));
   NOR2_X1 i_1_1_1073 (.A1(n_1_1_1156), .A2(n_1_1_1117), .ZN(n_1_1_1057));
   NOR2_X1 i_1_1_1074 (.A1(n_1_1_1159), .A2(n_1_1_1124), .ZN(n_1_1_1058));
   NOR2_X1 i_1_1_1075 (.A1(n_1_1_1172), .A2(n_1_1_1117), .ZN(n_1_1_1059));
   NOR2_X1 i_1_1_1076 (.A1(n_1_1_1154), .A2(n_1_1_1089), .ZN(n_1_1_1060));
   NOR2_X1 i_1_1_1077 (.A1(n_1_1_1136), .A2(n_1_1_1112), .ZN(n_1_1_1061));
   NOR2_X1 i_1_1_1078 (.A1(n_1_1_1176), .A2(n_1_1_1159), .ZN(n_1_1_1062));
   NOR2_X1 i_1_1_1079 (.A1(n_1_1_1112), .A2(n_1_1_1076), .ZN(n_1_1_1063));
   NOR2_X1 i_1_1_1080 (.A1(n_1_1_1169), .A2(n_1_1_1089), .ZN(n_1_1_1064));
   AOI22_X1 i_1_1_1081 (.A1(\mem[63] [15]), .A2(n_1_1_1116), .B1(n_1_1_1074), 
      .B2(\mem[9] [15]), .ZN(n_1_1_1065));
   NOR3_X1 i_1_1_1082 (.A1(n_1_1_1180), .A2(n_1_1_1164), .A3(n_1_1_1076), 
      .ZN(n_1));
   NOR2_X1 i_1_1_1083 (.A1(n_1_1_1164), .A2(n_1_1_1076), .ZN(n_1_1_1066));
   NOR3_X1 i_1_1_1084 (.A1(n_1_1_1180), .A2(n_1_1_1166), .A3(n_1_1_1076), 
      .ZN(n_2));
   NOR2_X1 i_1_1_1085 (.A1(n_1_1_1166), .A2(n_1_1_1076), .ZN(n_1_1_1067));
   NOR3_X1 i_1_1_1086 (.A1(n_1_1_1180), .A2(n_1_1_1169), .A3(n_1_1_1076), 
      .ZN(n_3));
   NOR2_X1 i_1_1_1087 (.A1(n_1_1_1169), .A2(n_1_1_1076), .ZN(n_1_1_1068));
   NOR3_X1 i_1_1_1088 (.A1(n_1_1_1180), .A2(n_1_1_1172), .A3(n_1_1_1076), 
      .ZN(n_4));
   NOR2_X1 i_1_1_1089 (.A1(n_1_1_1172), .A2(n_1_1_1076), .ZN(n_1_1_1069));
   NOR3_X1 i_1_1_1090 (.A1(n_1_1_1180), .A2(n_1_1_1176), .A3(n_1_1_1076), 
      .ZN(n_5));
   NOR2_X1 i_1_1_1091 (.A1(n_1_1_1176), .A2(n_1_1_1076), .ZN(n_1_1_1070));
   NOR3_X1 i_1_1_1092 (.A1(n_1_1_1180), .A2(n_1_1_1124), .A3(n_1_1_1076), 
      .ZN(n_6));
   NOR2_X1 i_1_1_1093 (.A1(n_1_1_1124), .A2(n_1_1_1076), .ZN(n_1_1_1071));
   NOR3_X1 i_1_1_1094 (.A1(n_1_1_1180), .A2(n_1_1_1143), .A3(n_1_1_1076), 
      .ZN(n_7));
   NOR2_X1 i_1_1_1095 (.A1(n_1_1_1143), .A2(n_1_1_1076), .ZN(n_1_1_1072));
   NOR2_X1 i_1_1_1096 (.A1(n_1_1_1098), .A2(n_1_1_1086), .ZN(n_8));
   NOR3_X1 i_1_1_1097 (.A1(n_1_1_1180), .A2(n_1_1_1128), .A3(n_1_1_1076), 
      .ZN(n_9));
   NOR2_X1 i_1_1_1098 (.A1(n_1_1_1128), .A2(n_1_1_1076), .ZN(n_1_1_1073));
   NOR3_X1 i_1_1_1099 (.A1(n_1_1_1180), .A2(n_1_1_1149), .A3(n_1_1_1076), 
      .ZN(n_10));
   NOR2_X1 i_1_1_1100 (.A1(n_1_1_1149), .A2(n_1_1_1076), .ZN(n_1_1_1074));
   NOR2_X1 i_1_1_1101 (.A1(n_1_1_1130), .A2(n_1_1_1085), .ZN(n_11));
   NOR2_X1 i_1_1_1102 (.A1(n_1_1_1130), .A2(n_1_1_1086), .ZN(n_12));
   NOR2_X1 i_1_1_1103 (.A1(n_1_1_1132), .A2(n_1_1_1085), .ZN(n_13));
   NOR3_X1 i_1_1_1104 (.A1(n_1_1_1180), .A2(n_1_1_1156), .A3(n_1_1_1076), 
      .ZN(n_14));
   NOR2_X1 i_1_1_1105 (.A1(n_1_1_1156), .A2(n_1_1_1076), .ZN(n_1_1_1075));
   NAND2_X1 i_1_1_1106 (.A1(n_1_1_1090), .A2(n_1_1_1187), .ZN(n_1_1_1076));
   NOR2_X1 i_1_1_1107 (.A1(n_1_1_1085), .A2(n_1_1_1077), .ZN(n_15));
   NOR2_X1 i_1_1_1108 (.A1(n_1_1_1086), .A2(n_1_1_1077), .ZN(n_16));
   NAND2_X1 i_1_1_1109 (.A1(n_1_1_1161), .A2(n_1_1_1131), .ZN(n_1_1_1077));
   NOR3_X1 i_1_1_1110 (.A1(n_1_1_1180), .A2(n_1_1_1164), .A3(n_1_1_1089), 
      .ZN(n_17));
   NOR2_X1 i_1_1_1111 (.A1(n_1_1_1164), .A2(n_1_1_1089), .ZN(n_1_1_1078));
   NOR2_X1 i_1_1_1112 (.A1(n_1_1_1086), .A2(n_1_1_1079), .ZN(n_18));
   NAND2_X1 i_1_1_1113 (.A1(n_1_1_1173), .A2(n_1_1_1147), .ZN(n_1_1_1079));
   NOR2_X1 i_1_1_1114 (.A1(n_1_1_1140), .A2(n_1_1_1085), .ZN(n_19));
   NOR3_X1 i_1_1_1115 (.A1(n_1_1_1180), .A2(n_1_1_1172), .A3(n_1_1_1089), 
      .ZN(n_20));
   NOR2_X1 i_1_1_1116 (.A1(n_1_1_1172), .A2(n_1_1_1089), .ZN(n_1_1_1080));
   NOR2_X1 i_1_1_1117 (.A1(n_1_1_1141), .A2(n_1_1_1085), .ZN(n_21));
   NOR3_X1 i_1_1_1118 (.A1(n_1_1_1180), .A2(n_1_1_1124), .A3(n_1_1_1089), 
      .ZN(n_22));
   NOR2_X1 i_1_1_1119 (.A1(n_1_1_1124), .A2(n_1_1_1089), .ZN(n_1_1_1081));
   NOR2_X1 i_1_1_1120 (.A1(n_1_1_1085), .A2(n_1_1_1082), .ZN(n_23));
   NOR2_X1 i_1_1_1121 (.A1(n_1_1_1086), .A2(n_1_1_1082), .ZN(n_24));
   NAND3_X1 i_1_1_1122 (.A1(address[4]), .A2(address[1]), .A3(n_1_1_1178), 
      .ZN(n_1_1_1082));
   NOR3_X1 i_1_1_1123 (.A1(n_1_1_1180), .A2(n_1_1_1128), .A3(n_1_1_1089), 
      .ZN(n_25));
   NOR2_X1 i_1_1_1124 (.A1(n_1_1_1128), .A2(n_1_1_1089), .ZN(n_1_1_1083));
   NOR3_X1 i_1_1_1125 (.A1(n_1_1_1180), .A2(n_1_1_1149), .A3(n_1_1_1089), 
      .ZN(n_26));
   NOR2_X1 i_1_1_1126 (.A1(n_1_1_1149), .A2(n_1_1_1089), .ZN(n_1_1_1084));
   NOR2_X1 i_1_1_1127 (.A1(n_1_1_1151), .A2(n_1_1_1085), .ZN(n_27));
   NOR2_X1 i_1_1_1128 (.A1(n_1_1_1151), .A2(n_1_1_1086), .ZN(n_28));
   NOR2_X1 i_1_1_1129 (.A1(n_1_1_1114), .A2(n_1_1_1085), .ZN(n_29));
   NAND3_X1 i_1_1_1130 (.A1(n_1_1_1179), .A2(n_1_1_1090), .A3(n_1_1_1184), 
      .ZN(n_1_1_1085));
   NOR2_X1 i_1_1_1131 (.A1(n_1_1_1114), .A2(n_1_1_1086), .ZN(n_30));
   NAND3_X1 i_1_1_1132 (.A1(address[0]), .A2(n_1_1_1179), .A3(n_1_1_1090), 
      .ZN(n_1_1_1086));
   NOR3_X1 i_1_1_1133 (.A1(n_1_1_1180), .A2(n_1_1_1158), .A3(n_1_1_1089), 
      .ZN(n_31));
   NOR2_X1 i_1_1_1134 (.A1(n_1_1_1158), .A2(n_1_1_1089), .ZN(n_1_1_1087));
   NOR3_X1 i_1_1_1135 (.A1(n_1_1_1180), .A2(n_1_1_1137), .A3(n_1_1_1089), 
      .ZN(n_32));
   NOR2_X1 i_1_1_1136 (.A1(n_1_1_1137), .A2(n_1_1_1089), .ZN(n_1_1_1088));
   NAND2_X1 i_1_1_1137 (.A1(address[4]), .A2(n_1_1_1090), .ZN(n_1_1_1089));
   NOR2_X1 i_1_1_1138 (.A1(address[6]), .A2(address[5]), .ZN(n_1_1_1090));
   NOR3_X1 i_1_1_1139 (.A1(n_1_1_1180), .A2(n_1_1_1164), .A3(n_1_1_1103), 
      .ZN(n_33));
   NOR2_X1 i_1_1_1140 (.A1(n_1_1_1164), .A2(n_1_1_1103), .ZN(n_1_1_1091));
   NOR3_X1 i_1_1_1141 (.A1(n_1_1_1180), .A2(n_1_1_1166), .A3(n_1_1_1103), 
      .ZN(n_34));
   NOR2_X1 i_1_1_1142 (.A1(n_1_1_1166), .A2(n_1_1_1103), .ZN(n_1_1_1092));
   NOR3_X1 i_1_1_1143 (.A1(n_1_1_1180), .A2(n_1_1_1169), .A3(n_1_1_1103), 
      .ZN(n_35));
   NOR2_X1 i_1_1_1144 (.A1(n_1_1_1169), .A2(n_1_1_1103), .ZN(n_1_1_1093));
   NOR3_X1 i_1_1_1145 (.A1(n_1_1_1180), .A2(n_1_1_1172), .A3(n_1_1_1103), 
      .ZN(n_36));
   NOR2_X1 i_1_1_1146 (.A1(n_1_1_1172), .A2(n_1_1_1103), .ZN(n_1_1_1094));
   NOR3_X1 i_1_1_1147 (.A1(n_1_1_1180), .A2(n_1_1_1176), .A3(n_1_1_1103), 
      .ZN(n_37));
   NOR2_X1 i_1_1_1148 (.A1(n_1_1_1176), .A2(n_1_1_1103), .ZN(n_1_1_1095));
   NOR3_X1 i_1_1_1149 (.A1(n_1_1_1180), .A2(n_1_1_1124), .A3(n_1_1_1103), 
      .ZN(n_38));
   NOR2_X1 i_1_1_1150 (.A1(n_1_1_1124), .A2(n_1_1_1103), .ZN(n_1_1_1096));
   NOR3_X1 i_1_1_1151 (.A1(n_1_1_1180), .A2(n_1_1_1143), .A3(n_1_1_1103), 
      .ZN(n_39));
   NOR2_X1 i_1_1_1152 (.A1(n_1_1_1143), .A2(n_1_1_1103), .ZN(n_1_1_1097));
   NOR2_X1 i_1_1_1153 (.A1(n_1_1_1113), .A2(n_1_1_1098), .ZN(n_40));
   NAND2_X1 i_1_1_1154 (.A1(n_1_1_1178), .A2(n_1_1_1131), .ZN(n_1_1_1098));
   NOR3_X1 i_1_1_1155 (.A1(n_1_1_1180), .A2(n_1_1_1128), .A3(n_1_1_1103), 
      .ZN(n_41));
   NOR2_X1 i_1_1_1156 (.A1(n_1_1_1128), .A2(n_1_1_1103), .ZN(n_1_1_1099));
   NOR3_X1 i_1_1_1157 (.A1(n_1_1_1180), .A2(n_1_1_1149), .A3(n_1_1_1103), 
      .ZN(n_42));
   NOR2_X1 i_1_1_1158 (.A1(n_1_1_1149), .A2(n_1_1_1103), .ZN(n_1_1_1100));
   NOR2_X1 i_1_1_1159 (.A1(n_1_1_1130), .A2(n_1_1_1115), .ZN(n_43));
   NOR2_X1 i_1_1_1160 (.A1(n_1_1_1130), .A2(n_1_1_1113), .ZN(n_44));
   NOR2_X1 i_1_1_1161 (.A1(n_1_1_1132), .A2(n_1_1_1115), .ZN(n_45));
   NOR2_X1 i_1_1_1162 (.A1(n_1_1_1132), .A2(n_1_1_1113), .ZN(n_46));
   NOR3_X1 i_1_1_1163 (.A1(n_1_1_1180), .A2(n_1_1_1158), .A3(n_1_1_1103), 
      .ZN(n_47));
   NOR2_X1 i_1_1_1164 (.A1(n_1_1_1158), .A2(n_1_1_1103), .ZN(n_1_1_1101));
   NOR3_X1 i_1_1_1165 (.A1(n_1_1_1180), .A2(n_1_1_1137), .A3(n_1_1_1103), 
      .ZN(n_48));
   NOR2_X1 i_1_1_1166 (.A1(n_1_1_1137), .A2(n_1_1_1103), .ZN(n_1_1_1102));
   NAND3_X1 i_1_1_1167 (.A1(n_1_1_1189), .A2(n_1_1_1187), .A3(address[5]), 
      .ZN(n_1_1_1103));
   NOR3_X1 i_1_1_1168 (.A1(n_1_1_1180), .A2(n_1_1_1164), .A3(n_1_1_1117), 
      .ZN(n_49));
   NOR2_X1 i_1_1_1169 (.A1(n_1_1_1164), .A2(n_1_1_1117), .ZN(n_1_1_1104));
   NOR3_X1 i_1_1_1170 (.A1(n_1_1_1180), .A2(n_1_1_1166), .A3(n_1_1_1117), 
      .ZN(n_50));
   NOR2_X1 i_1_1_1171 (.A1(n_1_1_1166), .A2(n_1_1_1117), .ZN(n_1_1_1105));
   NOR2_X1 i_1_1_1172 (.A1(n_1_1_1140), .A2(n_1_1_1115), .ZN(n_51));
   NOR2_X1 i_1_1_1173 (.A1(n_1_1_1140), .A2(n_1_1_1113), .ZN(n_52));
   NOR2_X1 i_1_1_1174 (.A1(n_1_1_1141), .A2(n_1_1_1115), .ZN(n_53));
   NOR2_X1 i_1_1_1175 (.A1(n_1_1_1141), .A2(n_1_1_1113), .ZN(n_54));
   NOR3_X1 i_1_1_1176 (.A1(n_1_1_1180), .A2(n_1_1_1143), .A3(n_1_1_1117), 
      .ZN(n_55));
   NOR2_X1 i_1_1_1177 (.A1(n_1_1_1143), .A2(n_1_1_1117), .ZN(n_1_1_1106));
   NOR3_X1 i_1_1_1178 (.A1(n_1_1_1180), .A2(n_1_1_1145), .A3(n_1_1_1117), 
      .ZN(n_56));
   NOR2_X1 i_1_1_1179 (.A1(n_1_1_1145), .A2(n_1_1_1117), .ZN(n_1_1_1107));
   NOR2_X1 i_1_1_1180 (.A1(n_1_1_1146), .A2(n_1_1_1115), .ZN(n_57));
   NOR3_X1 i_1_1_1181 (.A1(n_1_1_1180), .A2(n_1_1_1149), .A3(n_1_1_1117), 
      .ZN(n_58));
   NOR2_X1 i_1_1_1182 (.A1(n_1_1_1149), .A2(n_1_1_1117), .ZN(n_1_1_1108));
   NOR3_X1 i_1_1_1183 (.A1(n_1_1_1180), .A2(n_1_1_1117), .A3(n_1_1_1110), 
      .ZN(n_59));
   NOR2_X1 i_1_1_1184 (.A1(n_1_1_1117), .A2(n_1_1_1110), .ZN(n_1_1_1109));
   NAND2_X1 i_1_1_1185 (.A1(n_1_1_1170), .A2(n_1_1_1152), .ZN(n_1_1_1110));
   NOR3_X1 i_1_1_1186 (.A1(n_1_1_1180), .A2(n_1_1_1117), .A3(n_1_1_1112), 
      .ZN(n_60));
   NOR2_X1 i_1_1_1187 (.A1(n_1_1_1117), .A2(n_1_1_1112), .ZN(n_1_1_1111));
   NAND3_X1 i_1_1_1188 (.A1(address[1]), .A2(address[0]), .A3(n_1_1_1152), 
      .ZN(n_1_1_1112));
   NOR2_X1 i_1_1_1189 (.A1(n_1_1_1115), .A2(n_1_1_1114), .ZN(n_61));
   NOR2_X1 i_1_1_1190 (.A1(n_1_1_1114), .A2(n_1_1_1113), .ZN(n_62));
   NAND4_X1 i_1_1_1191 (.A1(address[5]), .A2(address[0]), .A3(n_1_1_1179), 
      .A4(n_1_1_1189), .ZN(n_1_1_1113));
   NAND2_X1 i_1_1_1192 (.A1(n_1_1_1161), .A2(n_1_1_1147), .ZN(n_1_1_1114));
   NOR2_X1 i_1_1_1193 (.A1(n_1_1_1160), .A2(n_1_1_1115), .ZN(n_63));
   NAND4_X1 i_1_1_1194 (.A1(address[5]), .A2(n_1_1_1179), .A3(n_1_1_1184), 
      .A4(n_1_1_1189), .ZN(n_1_1_1115));
   NOR3_X1 i_1_1_1195 (.A1(n_1_1_1180), .A2(n_1_1_1137), .A3(n_1_1_1117), 
      .ZN(n_64));
   NOR2_X1 i_1_1_1196 (.A1(n_1_1_1137), .A2(n_1_1_1117), .ZN(n_1_1_1116));
   NAND3_X1 i_1_1_1197 (.A1(n_1_1_1189), .A2(address[5]), .A3(address[4]), 
      .ZN(n_1_1_1117));
   NOR3_X1 i_1_1_1198 (.A1(n_1_1_1180), .A2(n_1_1_1164), .A3(n_1_1_1136), 
      .ZN(n_65));
   NOR2_X1 i_1_1_1199 (.A1(n_1_1_1164), .A2(n_1_1_1136), .ZN(n_1_1_1118));
   NOR3_X1 i_1_1_1200 (.A1(n_1_1_1180), .A2(n_1_1_1166), .A3(n_1_1_1136), 
      .ZN(n_66));
   NOR2_X1 i_1_1_1201 (.A1(n_1_1_1166), .A2(n_1_1_1136), .ZN(n_1_1_1119));
   NOR3_X1 i_1_1_1202 (.A1(n_1_1_1180), .A2(n_1_1_1169), .A3(n_1_1_1136), 
      .ZN(n_67));
   NOR2_X1 i_1_1_1203 (.A1(n_1_1_1169), .A2(n_1_1_1136), .ZN(n_1_1_1120));
   NOR3_X1 i_1_1_1204 (.A1(n_1_1_1180), .A2(n_1_1_1172), .A3(n_1_1_1136), 
      .ZN(n_68));
   NOR2_X1 i_1_1_1205 (.A1(n_1_1_1172), .A2(n_1_1_1136), .ZN(n_1_1_1121));
   NOR3_X1 i_1_1_1206 (.A1(n_1_1_1180), .A2(n_1_1_1176), .A3(n_1_1_1136), 
      .ZN(n_69));
   NOR2_X1 i_1_1_1207 (.A1(n_1_1_1176), .A2(n_1_1_1136), .ZN(n_1_1_1122));
   NOR3_X1 i_1_1_1208 (.A1(n_1_1_1180), .A2(n_1_1_1136), .A3(n_1_1_1124), 
      .ZN(n_70));
   NOR2_X1 i_1_1_1209 (.A1(n_1_1_1136), .A2(n_1_1_1124), .ZN(n_1_1_1123));
   NAND2_X1 i_1_1_1210 (.A1(n_1_1_1178), .A2(n_1_1_1167), .ZN(n_1_1_1124));
   NOR3_X1 i_1_1_1211 (.A1(n_1_1_1180), .A2(n_1_1_1143), .A3(n_1_1_1136), 
      .ZN(n_71));
   NOR2_X1 i_1_1_1212 (.A1(n_1_1_1143), .A2(n_1_1_1136), .ZN(n_1_1_1125));
   NOR3_X1 i_1_1_1213 (.A1(n_1_1_1180), .A2(n_1_1_1145), .A3(n_1_1_1136), 
      .ZN(n_72));
   NOR2_X1 i_1_1_1214 (.A1(n_1_1_1145), .A2(n_1_1_1136), .ZN(n_1_1_1126));
   NOR3_X1 i_1_1_1215 (.A1(n_1_1_1180), .A2(n_1_1_1136), .A3(n_1_1_1128), 
      .ZN(n_73));
   NOR2_X1 i_1_1_1216 (.A1(n_1_1_1136), .A2(n_1_1_1128), .ZN(n_1_1_1127));
   NAND2_X1 i_1_1_1217 (.A1(n_1_1_1177), .A2(n_1_1_1152), .ZN(n_1_1_1128));
   NOR3_X1 i_1_1_1218 (.A1(n_1_1_1180), .A2(n_1_1_1149), .A3(n_1_1_1136), 
      .ZN(n_74));
   NOR2_X1 i_1_1_1219 (.A1(n_1_1_1149), .A2(n_1_1_1136), .ZN(n_1_1_1129));
   NOR2_X1 i_1_1_1220 (.A1(n_1_1_1150), .A2(n_1_1_1130), .ZN(n_75));
   NOR2_X1 i_1_1_1221 (.A1(n_1_1_1162), .A2(n_1_1_1130), .ZN(n_76));
   NAND2_X1 i_1_1_1222 (.A1(n_1_1_1152), .A2(n_1_1_1131), .ZN(n_1_1_1130));
   NOR2_X1 i_1_1_1223 (.A1(n_1_1_1185), .A2(address[4]), .ZN(n_1_1_1131));
   NOR2_X1 i_1_1_1224 (.A1(n_1_1_1150), .A2(n_1_1_1132), .ZN(n_77));
   NAND3_X1 i_1_1_1225 (.A1(n_1_1_1161), .A2(n_1_1_1185), .A3(n_1_1_1187), 
      .ZN(n_1_1_1132));
   NOR3_X1 i_1_1_1226 (.A1(n_1_1_1180), .A2(n_1_1_1156), .A3(n_1_1_1136), 
      .ZN(n_78));
   NOR2_X1 i_1_1_1227 (.A1(n_1_1_1156), .A2(n_1_1_1136), .ZN(n_1_1_1133));
   NOR3_X1 i_1_1_1228 (.A1(n_1_1_1180), .A2(n_1_1_1158), .A3(n_1_1_1136), 
      .ZN(n_79));
   NOR2_X1 i_1_1_1229 (.A1(n_1_1_1158), .A2(n_1_1_1136), .ZN(n_1_1_1134));
   NOR3_X1 i_1_1_1230 (.A1(n_1_1_1180), .A2(n_1_1_1137), .A3(n_1_1_1136), 
      .ZN(n_80));
   NOR2_X1 i_1_1_1231 (.A1(n_1_1_1137), .A2(n_1_1_1136), .ZN(n_1_1_1135));
   NAND3_X1 i_1_1_1232 (.A1(n_1_1_1188), .A2(n_1_1_1187), .A3(address[6]), 
      .ZN(n_1_1_1136));
   NAND3_X1 i_1_1_1233 (.A1(address[1]), .A2(address[0]), .A3(n_1_1_1161), 
      .ZN(n_1_1_1137));
   NOR3_X1 i_1_1_1234 (.A1(n_1_1_1180), .A2(n_1_1_1164), .A3(n_1_1_1159), 
      .ZN(n_81));
   NOR2_X1 i_1_1_1235 (.A1(n_1_1_1164), .A2(n_1_1_1159), .ZN(n_1_1_1138));
   NOR3_X1 i_1_1_1236 (.A1(n_1_1_1180), .A2(n_1_1_1166), .A3(n_1_1_1159), 
      .ZN(n_82));
   NOR2_X1 i_1_1_1237 (.A1(n_1_1_1166), .A2(n_1_1_1159), .ZN(n_1_1_1139));
   NOR2_X1 i_1_1_1238 (.A1(n_1_1_1150), .A2(n_1_1_1140), .ZN(n_83));
   NOR2_X1 i_1_1_1239 (.A1(n_1_1_1162), .A2(n_1_1_1140), .ZN(n_84));
   NAND3_X1 i_1_1_1240 (.A1(address[4]), .A2(address[1]), .A3(n_1_1_1173), 
      .ZN(n_1_1_1140));
   NOR2_X1 i_1_1_1241 (.A1(n_1_1_1150), .A2(n_1_1_1141), .ZN(n_85));
   NOR2_X1 i_1_1_1242 (.A1(n_1_1_1162), .A2(n_1_1_1141), .ZN(n_86));
   NAND2_X1 i_1_1_1243 (.A1(n_1_1_1178), .A2(n_1_1_1147), .ZN(n_1_1_1141));
   NOR3_X1 i_1_1_1244 (.A1(n_1_1_1180), .A2(n_1_1_1159), .A3(n_1_1_1143), 
      .ZN(n_87));
   NOR2_X1 i_1_1_1245 (.A1(n_1_1_1159), .A2(n_1_1_1143), .ZN(n_1_1_1142));
   NAND2_X1 i_1_1_1246 (.A1(n_1_1_1178), .A2(n_1_1_1170), .ZN(n_1_1_1143));
   NOR3_X1 i_1_1_1247 (.A1(n_1_1_1180), .A2(n_1_1_1159), .A3(n_1_1_1145), 
      .ZN(n_88));
   NOR2_X1 i_1_1_1248 (.A1(n_1_1_1159), .A2(n_1_1_1145), .ZN(n_1_1_1144));
   NAND3_X1 i_1_1_1249 (.A1(address[1]), .A2(address[0]), .A3(n_1_1_1178), 
      .ZN(n_1_1_1145));
   NOR2_X1 i_1_1_1250 (.A1(n_1_1_1150), .A2(n_1_1_1146), .ZN(n_89));
   NAND2_X1 i_1_1_1251 (.A1(n_1_1_1152), .A2(n_1_1_1147), .ZN(n_1_1_1146));
   NOR2_X1 i_1_1_1252 (.A1(n_1_1_1187), .A2(address[1]), .ZN(n_1_1_1147));
   NOR3_X1 i_1_1_1253 (.A1(n_1_1_1180), .A2(n_1_1_1159), .A3(n_1_1_1149), 
      .ZN(n_90));
   NOR2_X1 i_1_1_1254 (.A1(n_1_1_1159), .A2(n_1_1_1149), .ZN(n_1_1_1148));
   NAND2_X1 i_1_1_1255 (.A1(n_1_1_1167), .A2(n_1_1_1152), .ZN(n_1_1_1149));
   NOR2_X1 i_1_1_1256 (.A1(n_1_1_1151), .A2(n_1_1_1150), .ZN(n_91));
   NAND4_X1 i_1_1_1257 (.A1(n_1_1_1188), .A2(n_1_1_1179), .A3(n_1_1_1184), 
      .A4(address[6]), .ZN(n_1_1_1150));
   NOR2_X1 i_1_1_1258 (.A1(n_1_1_1162), .A2(n_1_1_1151), .ZN(n_92));
   NAND3_X1 i_1_1_1259 (.A1(address[4]), .A2(address[1]), .A3(n_1_1_1152), 
      .ZN(n_1_1_1151));
   AND2_X1 i_1_1_1260 (.A1(n_1_1_1186), .A2(address[3]), .ZN(n_1_1_1152));
   NOR3_X1 i_1_1_1261 (.A1(n_1_1_1180), .A2(n_1_1_1159), .A3(n_1_1_1154), 
      .ZN(n_93));
   NOR2_X1 i_1_1_1262 (.A1(n_1_1_1159), .A2(n_1_1_1154), .ZN(n_1_1_1153));
   NAND2_X1 i_1_1_1263 (.A1(n_1_1_1177), .A2(n_1_1_1161), .ZN(n_1_1_1154));
   NOR3_X1 i_1_1_1264 (.A1(n_1_1_1180), .A2(n_1_1_1159), .A3(n_1_1_1156), 
      .ZN(n_94));
   NOR2_X1 i_1_1_1265 (.A1(n_1_1_1159), .A2(n_1_1_1156), .ZN(n_1_1_1155));
   NAND2_X1 i_1_1_1266 (.A1(n_1_1_1167), .A2(n_1_1_1161), .ZN(n_1_1_1156));
   NOR3_X1 i_1_1_1267 (.A1(n_1_1_1180), .A2(n_1_1_1159), .A3(n_1_1_1158), 
      .ZN(n_95));
   NOR2_X1 i_1_1_1268 (.A1(n_1_1_1159), .A2(n_1_1_1158), .ZN(n_1_1_1157));
   NAND2_X1 i_1_1_1269 (.A1(n_1_1_1170), .A2(n_1_1_1161), .ZN(n_1_1_1158));
   NAND3_X1 i_1_1_1270 (.A1(n_1_1_1188), .A2(address[4]), .A3(address[6]), 
      .ZN(n_1_1_1159));
   NOR2_X1 i_1_1_1271 (.A1(n_1_1_1162), .A2(n_1_1_1160), .ZN(n_96));
   NAND3_X1 i_1_1_1272 (.A1(address[4]), .A2(address[1]), .A3(n_1_1_1161), 
      .ZN(n_1_1_1160));
   AND2_X1 i_1_1_1273 (.A1(address[3]), .A2(address[2]), .ZN(n_1_1_1161));
   NAND4_X1 i_1_1_1274 (.A1(address[6]), .A2(n_1_1_1179), .A3(n_1_1_1188), 
      .A4(address[0]), .ZN(n_1_1_1162));
   NOR3_X1 i_1_1_1275 (.A1(n_1_1_1180), .A2(n_1_1_1175), .A3(n_1_1_1164), 
      .ZN(n_97));
   NOR2_X1 i_1_1_1276 (.A1(n_1_1_1175), .A2(n_1_1_1164), .ZN(n_1_1_1163));
   NAND2_X1 i_1_1_1277 (.A1(n_1_1_1177), .A2(n_1_1_1173), .ZN(n_1_1_1164));
   NOR3_X1 i_1_1_1278 (.A1(n_1_1_1180), .A2(n_1_1_1175), .A3(n_1_1_1166), 
      .ZN(n_98));
   NOR2_X1 i_1_1_1279 (.A1(n_1_1_1175), .A2(n_1_1_1166), .ZN(n_1_1_1165));
   NAND2_X1 i_1_1_1280 (.A1(n_1_1_1173), .A2(n_1_1_1167), .ZN(n_1_1_1166));
   NOR2_X1 i_1_1_1281 (.A1(n_1_1_1184), .A2(address[1]), .ZN(n_1_1_1167));
   NOR3_X1 i_1_1_1282 (.A1(n_1_1_1180), .A2(n_1_1_1175), .A3(n_1_1_1169), 
      .ZN(n_99));
   NOR2_X1 i_1_1_1283 (.A1(n_1_1_1175), .A2(n_1_1_1169), .ZN(n_1_1_1168));
   NAND2_X1 i_1_1_1284 (.A1(n_1_1_1173), .A2(n_1_1_1170), .ZN(n_1_1_1169));
   NOR2_X1 i_1_1_1285 (.A1(n_1_1_1185), .A2(address[0]), .ZN(n_1_1_1170));
   NOR3_X1 i_1_1_1286 (.A1(n_1_1_1180), .A2(n_1_1_1175), .A3(n_1_1_1172), 
      .ZN(n_100));
   NOR2_X1 i_1_1_1287 (.A1(n_1_1_1175), .A2(n_1_1_1172), .ZN(n_1_1_1171));
   NAND3_X1 i_1_1_1288 (.A1(address[1]), .A2(address[0]), .A3(n_1_1_1173), 
      .ZN(n_1_1_1172));
   NOR2_X1 i_1_1_1289 (.A1(address[3]), .A2(address[2]), .ZN(n_1_1_1173));
   NOR3_X1 i_1_1_1290 (.A1(n_1_1_1180), .A2(n_1_1_1176), .A3(n_1_1_1175), 
      .ZN(n_101));
   NOR2_X1 i_1_1_1291 (.A1(n_1_1_1176), .A2(n_1_1_1175), .ZN(n_1_1_1174));
   NAND3_X1 i_1_1_1292 (.A1(n_1_1_1187), .A2(address[5]), .A3(address[6]), 
      .ZN(n_1_1_1175));
   NAND2_X1 i_1_1_1293 (.A1(n_1_1_1178), .A2(n_1_1_1177), .ZN(n_1_1_1176));
   NOR2_X1 i_1_1_1294 (.A1(address[1]), .A2(address[0]), .ZN(n_1_1_1177));
   NOR2_X1 i_1_1_1295 (.A1(n_1_1_1186), .A2(address[3]), .ZN(n_1_1_1178));
   INV_X1 i_1_1_1296 (.A(n_1_1_1180), .ZN(n_1_1_1179));
   NAND3_X1 i_1_1_1297 (.A1(n_1_1_1183), .A2(n_1_1_1182), .A3(n_1_1_1181), 
      .ZN(n_1_1_1180));
   NOR4_X1 i_1_1_1298 (.A1(read_signal), .A2(n_1_1_1190), .A3(address[15]), 
      .A4(address[14]), .ZN(n_1_1_1181));
   NOR4_X1 i_1_1_1299 (.A1(address[13]), .A2(address[12]), .A3(address[11]), 
      .A4(address[10]), .ZN(n_1_1_1182));
   NOR3_X1 i_1_1_1300 (.A1(address[9]), .A2(address[8]), .A3(address[7]), 
      .ZN(n_1_1_1183));
   INV_X1 i_1_1_1301 (.A(address[0]), .ZN(n_1_1_1184));
   INV_X1 i_1_1_1302 (.A(address[1]), .ZN(n_1_1_1185));
   INV_X1 i_1_1_1303 (.A(address[2]), .ZN(n_1_1_1186));
   INV_X1 i_1_1_1304 (.A(address[4]), .ZN(n_1_1_1187));
   INV_X1 i_1_1_1305 (.A(address[5]), .ZN(n_1_1_1188));
   INV_X1 i_1_1_1306 (.A(address[6]), .ZN(n_1_1_1189));
   INV_X1 i_1_1_1307 (.A(write_signal), .ZN(n_1_1_1190));
endmodule
